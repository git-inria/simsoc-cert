Require Import Globalenvs Memory.
Require Import Csyntax Csem Cstrategy Coqlib Integers Values Maps Errors. 
Require Import Arm6_State Arm6_Proc Arm6_SCC Bitvec Arm6.
Require Import adc_compcert_fixed.
Require Import projection. 

Require Import Arm6_Simul.
Import I.
Import Arm6_Functions.Semantics.

(* Functional relation between the C memory module which contains the other ADC parameters, 
   and the COQ specification of ADC parameters *)
Definition sbit_func_related (m:Mem.mem) (e:env) (sbit:bool):Prop:=
  bit_proj m e S = sbit.

Definition cond_func_related (m:Mem.mem) (e:env) (cond:opcode):Prop:=
  cond_proj m e = cond.

Definition d_func_related (m:Mem.mem) (e:env) (d:regnum):Prop:=
  reg_proj m e adc_compcert_fixed.d = d.

Definition n_func_related (m:Mem.mem) (e:env) (n:regnum):Prop:=
  reg_proj m e adc_compcert_fixed.n = n.

Definition so_func_related (m:Mem.mem) (e:env) (so:word):Prop:=
  bits_proj m e shifter_operand = so.

(* Human readable renaming of [p], which is generated by the Coq printer *)
(*Definition prog_adc := adc_compcert_fixed.p.*)

(* The assignment of old_Rn has a normal outcome *)
Lemma normal_outcome_for_assgnt: 
  forall a1 a2 ge t ev m e m' out,
  exec_stmt ge e m (Sdo (Eassign a1 a2 t)) ev m' out ->
  out = Out_normal.
Proof.
intros until out. intros exst. 
inv exst. reflexivity.
Qed.

Implicit Arguments normal_outcome_for_assgnt [a1 a2 ge t ev m e m' out].

Ltac noa :=
  match goal with
    [He: exec_stmt _ _ _ (Sdo (Eassign _ _ _)) _ _ ?out,
     Hd: ?out <> Out_normal |- _ ] =>
       case Hd; 
       apply (normal_outcome_for_assgnt He) end.

(* Any Sdo has a normal outcome*)
Lemma normal_outcome_for_do:
  forall exp ge t m e m' out,
    exec_stmt ge e m (Sdo exp) t m' out ->
    out = Out_normal.
Proof.
  intros until out. intros exst.
  inv exst. reflexivity.
Qed.

Implicit Arguments normal_outcome_for_do [exp ge t m e m' out].

Ltac nod :=
  match goal with
    [He: exec_stmt _ _ _ (Sdo _) _ _ ?out,
     Hd: ?out <> Out_normal |- _ ] =>
       case Hd; 
       apply (normal_outcome_for_do He) end.  

(* Return the memory model which only relates to this ident *)
Parameter of_mem : AST.ident -> Mem.mem -> Mem.mem.

(*exp get_bit*)
Print fun_internal_ADC.

Definition reg_id id :=
  Ecall (Evalof (Evar reg T2) T2)
  (Econs (Evalof (Evar proc T3) T3)
    (Econs 
      (Evalof (Evar id T4) T4) Enil)) T1.

Definition get_rd_bit31 :=
  Ecall (Evalof (Evar get_bit T16) T16)
  (Econs (reg_id d)
    (Econs (Eval (Vint (repr 31)) T9)
      Enil)) T4.

Lemma same_reg_d :
  forall e m t m' a' l b st d,
    proc_state_related m e (Ok tt (mk_semstate l b st)) ->
    d_func_related m e d ->    
    eval_expr (Genv.globalenv prog_adc) e m RV 
              (reg_id adc_compcert_fixed.d) t m' a' ->
    a'= (Eval (Vint (Arm6_State.reg_content st d)) T1).
Admitted.

Set Implicit Arguments.

Lemma alloc_diff_block :
  forall m e e' m' x y b_x tx b_y ty,
    alloc_variables e m ((x,tx)::(y,ty)::nil) e' m'->
    list_norepet (x::y::nil) ->
    e' ! x = Some (b_x, tx) ->
    e' ! y = Some (b_y, ty) ->
    b_x <> b_y.
Proof.
  intros until ty. intros av norepet getx gety.
  inv av. inv H7. inv H9.
  apply Mem.valid_new_block in H6.
  unfold Mem.valid_block in H6.
  apply Mem.alloc_result in H8.
  rewrite <- H8 in H6; clear H8.
(* SearchPattern (_ < _ -> _ <> _). *)
  apply Zlt_not_eq in H6.
  assert (findy: (PTree.set y (b0, ty) (PTree.set x (b1, tx) e)) ! y =
                  Some (b0, ty)).
  apply PTree.gss. rewrite findy in gety. inversion gety.

  assert (findx: (PTree.set y (b0, ty) (PTree.set x (b1, tx) e)) ! x =
                  (PTree.set x (b1, tx) e) ! x).
  apply PTree.gso.
  inv norepet. unfold In in H2. intro exy. apply H2. left. symmetry. exact exy.

(*info intuition.*)

  rewrite findx in getx.
  rewrite PTree.gss in getx. inversion getx.
  rewrite <- H0. rewrite <- H1.
  exact H6.
Qed.

Set Printing Depth 30.
(*
Lemma and_zdiv_1:
  forall (x:word) (n:Z),
    0 < n < Z_of_nat wordsize ->
    (repr n) = x -> and (repr n) x / n = 1.
Proof.
  intros. rewrite <- H0. SearchAbout and. rewrite and_idem.
  SearchAbout Zdiv. 
*)
Lemma same_getbit :
  forall x n ,
    0 < n < Z_of_nat wordsize ->
    zero_ext 8 (and (shru x (repr n)) (repr 1)) = x [nat_of_Z n].
Proof.
  intros.
  assert (0 < 8 < Z_of_nat wordsize).
  simpl. omega.
  apply zero_ext_and with (x := (and (shru x (repr n)) (repr 1))) in H0.
  rewrite H0.  
  unfold bit. unfold bits. unfold bits_val.
  unfold masks. (*SearchAbout minus. *)
  rewrite minus_diag. (*Print masks_aux.*)
  simpl masks_aux. 
  (*SearchAbout repr.*)
  rewrite shru_div_two_p.

(*
  induction n. 
  simpl nat_of_Z. 
  unfold masks. simpl masks_aux.
  rewrite two_power_nat_O.
  SearchAbout (Zdiv).
  rewrite Zdiv_1_r.
  (*lemma on 'repr' apply eqm_samerepr. apply eqm_refl2.*)
  SearchAbout two_p.
  assert (8 = Z_of_nat 8).
  simpl; reflexivity. rewrite H0.
  rewrite <- two_power_nat_two_p.
  rewrite Word.shru_zero.
  SearchAbout and.
  admit.
  admit.
  unfold nat_of_Z.
  unfold masks. simpl masks_aux.
  rewrite two_power_nat_O.
  rewrite Zdiv_1_r.
  assert (8 = Z_of_nat 8).
  simpl; reflexivity. rewrite H0.
  rewrite <- two_power_nat_two_p.
  SearchAbout Zneg.
*)
Admitted.

(* expirement on how to avoid using inversion *)
(*
Ltac gen_inv_S y :=
 pattern y; 
 match goal with [ |- ?concl _ ] => 
   change (match S y with S y => concl y | _ => True end) end;
 cbv beta.
*)

Ltac case_I h := case h; try (intros; exact I); clear h.

Ltac case_h h := case h; clear h; try contradiction.

Ltac rew_clean eq :=
  match type of eq with ?l = ?r => rewrite eq in *; clear eq l end.

Ltac and_eq_subst ae :=
  repeat (rew_clean ae) ||
         (let feq := fresh "eq" in destruct ae as [feq ae];
          rew_clean feq).

Ltac inv_end ev mm mm' :=
   unfold ev, mm, mm' in *; clear ev mm mm'; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_ecall_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env arg_m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?c] =>
    pose (e := Ecall a1 a2 a3); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert 
      (em : match e with 
                      |Ecall a b c =>
                        (a=a1)/\(b=a2)/\(c=a3)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                      |_=> False
                    end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.

Ltac inv_ecall arg_m t1 m2 rf' t2 m3 rargs' 
         vf vargs0 targs tres fd t3 vres H H0 H1 H2 H3 H4 H5 H6 :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_ecall_begin arg_m ev mm mm'; 
  intros e0 m1 rf rargs ty t1 m2 rf' t2 m3 rargs' 
         vf vargs0 targs tres fd t3 m4 vres H H0 H1 H2 H3 H4 H5 H6;
  inv_end ev mm mm'.

Ltac inv_evalof_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env arg_m _ (Evalof ?a1 ?a2) _ ?m' _ |- ?c ] =>
    pose (e := Evalof a1 a2); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert 
      (em : match e with 
                    |Evalof a b => 
                      (a=a1)/\(b=a2)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                    |_ => False
                  end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.

Ltac inv_evalof arg_m t0 m'0 a' H :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_evalof_begin arg_m ev mm mm'; 
  intros e0 m1 a t0 m'0 a' ty H;
  inv_end ev mm mm'.

Ltac inv_evar_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h: eval_expr _ ?env arg_m _ (Evar ?a1 ?a2) _ ?m' _ |- ?c] =>
    pose (e := Evar a1 a2); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert
      (em: match e with
                   |Evar a b => 
                     (a=a1)/\(b=a2)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                   |_ => False
                 end)
      by repeat (split||reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.
  
Ltac inv_evar arg_m :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_evar_begin arg_m ev mm mm';
  intros e0 m1 x ty;
  inv_end ev mm mm'. 

Ltac inv_evalof_simplrv_begin v :=
  match goal with [h: eval_simple_rvalue _ _ _ (Evalof ?a1 ?a2) v |- ?c] =>
    let e := fresh "expr" in
    pose (e := Evalof a1 a2);
    assert
      (rm: match e with
                   |Evalof a b =>(a = a1) /\ (b = a2)
                   |_=>False
                 end)
      by repeat  (split||reflexivity);
    fold e in h;
    revert rm;
    case_h h;
    clear e
  end.

Ltac inv_evalof_simplrv_end :=
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_evalof_simplrv v b0 ofs v0 H H0 H1 :=
  inv_evalof_simplrv_begin v;
  intros b0 ofs l0 ty v0 H H0 H1;
  inv_evalof_simplrv_end. 

Ltac inv_av_cons_begin arg_m ev :=
  let lst := fresh "lst" in
  match goal with [av: alloc_variables ?env arg_m ((?id,?ty) ::?t) ?a3 ?a4 |- ?c] => 
    pose (lst := ((id,ty)::t)); pose (ev:=env);
    change (alloc_variables ev arg_m lst a3 a4) in av;
    assert
      (lm: match lst with
                    |(a,b)::c=>(a=id)/\(b=ty)/\(c=t)/\(ev=env)
                    |_=>False
                  end)
      by repeat (split||reflexivity);
    revert lm;
    case_h av;
    clear lst
  end.

Ltac inv_av_cons_end ev :=
   unfold ev in *; clear ev; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).  

Ltac inv_av_cons arg_m m m1 b1 m4 e2 H H0:=
  let ev:=fresh "ev" in 
  inv_av_cons_begin arg_m ev;
  intros e0 m id0 ty vars m1 b1 m4 e2 H H0;
  inv_av_cons_end ev.

Ltac inv_av_nil_begin arg_m lnil ev ev' :=  
  match goal with [av: alloc_variables ?env arg_m ?lst ?env' ?a4 |- ?c] =>
    pose (lnil:=lst); pose (ev:=env); pose (ev':=env');
    change (alloc_variables ev arg_m lnil ev' a4) in av;
    assert (lm:match lnil with 
                        |nil =>(nil = lst)/\(ev=env)/\(ev'=env')
                        |_ =>False end) 
      by repeat (split||reflexivity);
    revert lm;
    case_h av    
  end.

Ltac inv_av_nil_end lnil ev ev' :=
   unfold lnil, ev, ev' in *; clear lnil ev ev'; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_av_nil arg_m e0 m :=
  let lnil:=fresh "lnil" in 
  let ev:=fresh "ev" in 
  let ev':=fresh "ev'" in 
  inv_av_nil_begin arg_m lnil ev ev';
  intros e0 m;
  inv_av_nil_end lnil ev ev'.  

(*
Definition inv_expr_ecall e m ex m' (ex':expr):=
  match ex with
    |Ecall a b c => 
      forall (X:Prop), 
      (forall g t1 m1 rf' t2 m2 rargs' vf vargs targs tres fd t3 vres,
      eval_expr g e m RV a t1 m1 rf' -> 
      eval_exprlist g e m1 b t2 m2 rargs' ->
      eval_simple_rvalue g e m2 rf' vf ->
      eval_simple_list g e m2 rargs' targs vargs ->
      typeof a = Tfunction targs tres ->
      Genv.find_funct g vf = Some fd ->
      type_of_fundef fd = Tfunction targs tres ->
      eval_funcall g m2 fd vargs t3 m' vres -> X) -> X
    |_=> True
  end.
*)

Definition inv_expr_ecall' g e m ex m' ex':=
  match ex with
    |Ecall a b c =>
      forall (X:expr -> Prop),
      (forall t1 m1 rf' t2 m2 rargs' vf vargs targs tres fd t3 vres ty,
      eval_expr g e m RV a t1 m1 rf' -> 
      eval_exprlist g e m1 b t2 m2 rargs' ->
      eval_simple_rvalue g e m2 rf' vf ->
      eval_simple_list g e m2 rargs' targs vargs ->
      typeof a = Tfunction targs tres ->
      Genv.find_funct g vf = Some fd ->
      type_of_fundef fd = Tfunction targs tres ->
      eval_funcall g m2 fd vargs t3 m' vres -> 
      X (Eval vres ty)) -> X ex'
    |_=> True
  end.


Lemma same_get_reg' :
  forall e m0 m0' vargs m l b s d t m' v,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    proc_state_related m e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m get_rd_bit31  t m' v->
    v = Vint ((Arm6_State.reg_content s d) [n31]).
Proof.
  intros until v. intros av bp psrel dfrel get_bit.
  
  inversion get_bit as [env m1 gb t1 m1' gb' v1 gb_expr ev_rv Heqenv Heqm
    Heqexp Heqt Heqm' Heqv]; clear get_bit; subst.

  unfold get_rd_bit31 in gb_expr.

(*  revert ev_rv.
*)

(** new thought *)
(** Using impredicative encoding in inversion tactic *)
generalize 
  (match gb_expr in (eval_expr _ e m _ ex _ m' ex')
  return inv_expr_ecall' (Genv.globalenv prog_adc) e m ex m' ex' with
     |eval_call _ _ rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs
                      targs tres fd t3 _ vres H1 H2 H3 H4 H5 H6 H7 H8 =>
       (fun X k => k t1 m1 rf' t2 m2 rargs' vf vargs 
      targs tres fd t3 vres ty H1 H2 H3 H4 H5 H6 H7 H8 )
     |_=> I
   end). clear gb_expr.
intro k. red in k. revert ev_rv. apply k. clear k. 
intros until ty. 
intros gb_expr ev_explst ev_rv1 ev_simlst Heqty_gb Heqff Heqtyfd ev_funcall.
intro ev_rv.


(** Using impredicative encoding, 
   but without considering the output of expression evaluation *)
(*
generalize 
  (match gb_expr in (eval_expr _ e m _ ex _ m' ex')
  return inv_expr_ecall e m ex m' ex' with
     |eval_call e m rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs
                      targs tres fd t3 m3 vres H1 H2 H3 H4 H5 H6 H7 H8 =>
       (fun X k => k (Genv.globalenv prog_adc) t1 m1 rf' t2 m2 rargs' vf vargs 
                     targs tres fd t3 vres H1 H2 H3 H4 H5 H6 H7 H8)
     |_=> I
   end). clear gb_expr.
intro k. apply k. clear k.
*)

(** Without impredicative encoding *)
(* info 
  match goal with [h : eval_expr _ ?env ?m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?cl] =>
    let ex := fresh "expr_call" in
    pose (arg1 := a1);  
    pose (arg2 := a2);  
    pose (arg3 := a3);
    pose (ex := Ecall arg1 arg2 arg3);
    change (match ex with 
                      |Ecall a b c => cl
                      |_=> True
                    end);
    assert (ee : ex = Ecall arg1 arg2 arg3) by reflexivity; 
    revert ee;
    revert av bp psrel dfrel;
  
    change (Ecall a1 a2 a3) with ex in gb_expr;
    case gb_expr; try (intros; exact I); clear gb_expr e m t m' gb';
    intros e m rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs0 targs tres fd
      t3 m3 vres;
    intros gb_expr ev_exlst ev_simprv1 ev_simplst Heqtyrf Heqff Heqtyfd ev_funcall;
    intros av bp pstrl dfrel Heqexpr ev_simprv;
    injection Heqexpr; intros Heqty Heqrargs Heqrf;
    unfold arg1, arg2, arg3 in Heqty, Heqrargs, Heqrf; 
    clear arg1 arg2 arg3 Heqexpr expr_call;
    rewrite Heqty in ev_simprv;
    rewrite Heqrargs in ev_exlst;
    rewrite Heqrf in gb_expr, Heqtyrf;
    clear Heqty Heqrargs Heqrf
  end.
*)  

(* *********************************************************************)
(** old one *)
(** With extra equalities introduced in inversion tactic *)
(* 
Ltac inv_ecall_begin ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env ?m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?c] =>
    pose (e := Ecall a1 a2 a3); 
    pose (ev:=env); pose (mm:=m); pose (mm':=m');
    assert 
      (em : match e with 
                      |Ecall a b c =>
                        (a=a1)/\(b=a2)/\(c=a3)/\(env=ev)/\(m=mm)/\(m'=mm')
                      |_=> False
                    end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.
*)

(*
  inv_ecall m t1 m2 rf' t2 m3 rargs' vf vargs0 targs tres fd t3 vres
            gb_expr explst ev_rv1 ev_simlst H_ Heqfindfd Heqt16 ev_funcall. clear H_.
  intro ev_rv.
*)


(*
  (*harmless inversion: no ordering changes, no new hyp*)
  inversion ev_rv; subst; clear ev_rv.

  revert ev_rv1.
  inv_evalof m t0 m'0 a' H.
(*intro ev_rv1.

  revert ev_rv1.*)
  inv_evar m.
  intro ev_rv1.
  clear t0 a'.

  inv_evalof_simplrv vf b0 ofs v0 ev_simpl_lv Heqty Heqlvot.

  assert (globenv: e!get_bit=None).
    simpl in av.
    
    inv_av_cons m0 ma_proc m_proc b_proc m_proc' e_proc Heqma_proc av.
    inv_av_cons m_proc ma_s m_s b_s m_s' e_s Heqma_s av.
    inv_av_cons m_s ma_cond m_cond b_cond m_cond' e_cond Heqma_cond av.
    inv_av_cons m_cond ma_d m_d b_d m_d' e_d Heqma_d av.
    inv_av_cons m_d ma_n m_n b_n m_n' e_n Heqma_n av.
    inv_av_cons m_n ma_so m_so b_so m_so' e_so Heqma_so av.
    inv_av_cons m_so ma_on m_on b_on m_on' e_on Heqma_on av.

    inv_av_nil_begin m_on lnil ev ev'.
    intros.

    destruct lm as [feq ae]; clear feq.
    destruct ae as [feq ae]; rewrite feq in *; clear feq.
    rewrite <- ae in *; clear ae.

    
*)
    (*
    simpl; reflexivity.

  match goal with [_: eval_simple_lvalue _ _ _ (Evar ?a1 ?a2) _ _ |- ?c] =>
    assert
      (lv_match: match expr_evar with
                   |Evar a b =>(a = a1) /\ (b = a2)
                   |_=>False
                 end)
      by repeat  (split||reflexivity)
  end. 
  fold expr_evar in ev_lv.
  revert lv_match.

  case_h ev_lv.
    (*get_bit is in global environment *)
    intros until b1. intro locenv. intros.
    destruct lv_match as [eq1 eq2]; subst.
    rewrite locenv in globenv; discriminate.
    (*get_bit is in local environment *)
    intros until b1; intros _ Heqfindsymb _; intros.
    destruct lv_match as [eq1 eq2]; rewrite eq1 in *; clear eq1 eq2.*)

    (*match goal with [_:eval_exprlist _ _ _ (Econs ?a1 ?a2) _ _ _]*)
    
    
   
  

(* useful trick for later
  match goal with [_ : eval_expr _ _ _ _ ?interesting _ _ _ |- ?c ] => 
     let name := fresh e0 in 
     pose (name := interesting) end.
*)  

  (*revert gb_sim_rv.  
  generalize (refl_equal get_bit_reg).
  unfold get_bit_reg at 2.
  case gb_expr; clear gb_expr; try (intros; discriminate). 
  intros. injection H7. clear H7. intros; subst.*)


(*match goal with [ |- context c [Ecall ?a1 ?a2 ?a3]] => pattern a1, a2, a3 end.
    change 
      (match Ecall (Evalof (Evar get_bit T16) T16)
     (Econs (reg_id adc_compcert_fixed.d)
        (Econs (Eval (Vint (repr 31)) T9) Enil)) T4 with 
         | Ecall a b c => 
(fun (e0 : expr) (e1 : exprlist) (t0 : type) =>
    get_bit_reg = Ecall e0 e1 t0 ->
    v = Vint (Arm6_State.reg_content s d) [n31]) a b c
 | _ => True end). cbv beta.
  case_I gb_expr. red.
*)

(*
  generalize (refl_equal get_bit_reg).
  pattern get_bit_reg at 1.*)

  (*match goal with [ |- ?concl _ _ _ ] =>
    change 
      (match Ecall a1 a2 a3 with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  
  unfold get_bit_reg in gb_expr.
match goal with [ |- ?concl] => change ((fun _ _ _ => concl) 
   (Evalof (Evar get_bit T16) T16)
   (Econs (reg_id adc_compcert_fixed.d)
                    (Econs (Eval (Vint (repr 31)) T9) Enil))
   T4) end.
  match goal with [ gb_expr : context c [Ecall ?a1 ?a2 ?a3] |- ?concl _ _ _ ] =>
    change 
      (match Ecall a1 a2 a3 with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  case_I gb_expr. red.
  intros until rargs. intro ty.
  intros until vres.
  intros rf_exp rargs_exp vf_rval targs_vlst Heqtprf Heqfun Heqtpfun fd_funcall.
  
  match goal with [ |- ?concl _ _ _ ] =>
    change 
      (match get_bit_reg with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  

  case_eq get_bit_reg. intro
  case get_bit. intro
  unfold get_bit_reg in get_bit.*)
Admitted.



Lemma same_get_reg :
  forall e m0 m0' vargs m l b s d t m' v,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    proc_state_related m e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m get_rd_bit31 t m' v->
    v = Vint ((Arm6_State.reg_content s d) [n31]).
Proof.
  intros until v. intros av bp psrel dfrel get_bit.
  inv get_bit. 
  (*rename H into get_bit_reg_exp, H0 into get_bit_reg_v.
  inv get_bit_reg_exp.*) 
  inv H.
  inv H4. inv H8. inv H9. inv H5.
  
  (** HERE expand function reg *)



  apply same_reg_d with e m2 t1 m1 a1' l b s d in H4;
    [idtac| exact psrel |exact dfrel].
  rewrite H4 in *. 
  inv H13. inv H5. inv H14.
  inv H0. inv H6. inv H2. inv H4.

  assert (e!get_bit=None).
    inv av. inv H9. inv H13. inv H14. inv H15. inv H17. inv H18. inv H19.
    simpl. reflexivity.   
  assert (wdsz:0<31<Z_of_nat wordsize). unfold wordsize. unfold Wordsize_32.wordsize.
  simpl Z_of_nat. omega.
  inv H1.
    (*get_bit is in local env*)
    rewrite H in H5. discriminate H5.
    
    (*get_bit is in gloval env*)
    inv H7. inv H6. inv H13. inv H14. inv H6. simpl in H10, H9.
    inv H9.
    
      (*cast int to int*) 
      simpl in H16.
      inv H10; simpl in H16; inv H4; clear H8; inv H11;
        induction (eq_dec w0 w0);[idtac|inv H1|inv H4|inv H4].
      inv H1.
      clear H12.
      inv H16. inv H5. simpl in H6.
      destruct H6.
      inv H10. inv H6. inv H18. inv H17. inv H12. inv H20. inv H12. inv H19.
      inv H5; inv H7; simpl in H14; unfold sem_and in  H14; simpl in H14;
        [simpl|inv H9|inv H9].
      destruct v1,v2; inv H14. inv H13. inv H12. simpl in H14.
      inv H4. inv H19. inv H21. inv H11; clear H7. inv H13; clear H9.
      inv H6; [idtac| inv H11].
      inv H7; [idtac| inv H9].
      rewrite H13 in H17. rewrite H11 in H16.
      inv H17; inv H16.
      unfold load_value_of_type in *; simpl in H10, H12.
      unfold store_value_of_type in *; simpl in H18, H20.
      generalize H20; intro.
      apply Mem.load_store_other with
        AST.Mint32 _ _ _ _ _ AST.Mint32 b0 (signed w0) in H4.
      rewrite H4 in H10.
      eapply Mem.load_store_same in H20;[idtac|simpl; auto].
      rewrite H12 in H20.
      eapply Mem.load_store_same in H18;[idtac|simpl; auto].
      rewrite H10 in H18.
      inv H18; inv H20. inv H14.
      rewrite (same_getbit (Arm6_State.reg_content s d) wdsz). reflexivity.
      left. apply (alloc_diff_block H2); assumption.

      (*cast has no change*)
      clear H1; clear H2.
      clear H12.
      inv H16.
      inv H5. simpl in H6.
      destruct H6.
      inv H10. inv H6. inv H18. inv H17. inv H12. inv H20. inv H12. inv H19.
      inv H5; inv H7; simpl in H14; unfold sem_and in  H14; simpl in H14;
        [simpl|inv H9|inv H9].
      destruct v1,v2; inv H14. inv H13. inv H12. simpl in H14.
      inv H4. inv H19. inv H21. inv H11; clear H7. inv H13; clear H9.
      inv H6; [idtac| inv H11].
      inv H7; [idtac| inv H9].
      rewrite H13 in H17. rewrite H11 in H16.
      inv H17; inv H16.
      unfold load_value_of_type in *; simpl in H10, H12.
      unfold store_value_of_type in *; simpl in H18, H20.
      generalize H20; intro.
      apply Mem.load_store_other with
        AST.Mint32 _ _ _ _ _ AST.Mint32 b0 (signed w0) in H4.
      rewrite H4 in H10.
      eapply Mem.load_store_same in H20;[idtac|simpl; auto].
      rewrite H12 in H20.
      eapply Mem.load_store_same in H18;[idtac|simpl; auto].
      rewrite H10 in H18.
      inv H18; inv H20. inv H14.
      rewrite (same_getbit (Arm6_State.reg_content s d) wdsz); reflexivity.
      left. apply (alloc_diff_block H2); assumption.

      clear H1; clear H2.
      inv H4. inv H11; clear H8.
      induction (eq_dec w0 w0); [idtac|inv H1].
      inv H1. clear H12.
      inv H16.
      inv H5. simpl in H6. destruct H6.
      inv H5; [idtac|inv H7|inv H7].
      inv H11; inv H5; inv H19; inv H18; inv H17; inv H12; inv H19; inv H12.
      inv H4; inv H18; inv H20.
      inv H6. inv H12. inv H13. simpl in H14. simpl in H20.
      inv H11. inv H18.
      inv H7; inv H11.
      inv H6; [rewrite H13 in H16; inv H16|rewrite H7 in H16; inv H16].        
      inv H9; [rewrite H11 in H15; inv H15|rewrite H6 in H15; inv H15].
      unfold load_value_of_type in *; simpl in H12, H21.
      unfold store_value_of_type in *; simpl in H17, H19.
      inv H10; simpl in H17.

        (*cast int to int*)
        generalize H19; intro.
        apply Mem.load_store_other with
          AST.Mint32 _ _ _ _ _ AST.Mint32 b0 (signed w0) in H4.
        rewrite H4 in H12.
        eapply Mem.load_store_same in H17; [idtac|simpl; auto].
        simpl in H17.
        rewrite H17 in H12; inv H12.
        eapply Mem.load_store_same in H19; [idtac|simpl; auto].
        simpl in H19.
        rewrite H19 in H21; inv H21.
        unfold sem_shr in H20. simpl in H20. inv H20.
        inv H14. simpl.
        rewrite (same_getbit (Arm6_State.reg_content s d) wdsz); reflexivity.
        left. apply (alloc_diff_block H2); assumption.

        (*cast has no change*)
        generalize H19; intro.
        apply Mem.load_store_other with
          AST.Mint32 _ _ _ _ _ AST.Mint32 b0 (signed w0) in H4.
        rewrite H4 in H12.
        eapply Mem.load_store_same in H17; [idtac|simpl; auto].
        simpl in H17.
        rewrite H17 in H12; inv H12.
        eapply Mem.load_store_same in H19; [idtac|simpl; auto].
        simpl in H19.
        rewrite H19 in H21; inv H21.
        unfold sem_shr in H20. simpl in H20. inv H20.
        inv H14. simpl.
        rewrite (same_getbit (Arm6_State.reg_content s d) wdsz); reflexivity.
        left. apply (alloc_diff_block H2); assumption.
Qed.
          


Unset Implicit Arguments.
(* Assume that every function that ADC calls, executes correctly
   and the C proc and ARM state related after these function execution *)
Axiom functions_behavior_ok:
  forall e l b s vf fd m vargs t m' vres l' b' s',
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    Genv.find_funct (Genv.globalenv prog_adc) vf = Some fd ->
    eval_funcall (Genv.globalenv prog_adc) m fd vargs t m' vres ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l' b' s')).

(* Assume that call to unpredictable leads to an Ko result*)
Axiom funct_unpredictable:
  forall e semstt vf fd m vargs t m' vres,
    proc_state_related (of_mem proc m) e (Ok tt semstt) ->
    Genv.find_funct (Genv.globalenv prog_adc) vf = Some fd ->
    eval_funcall (Genv.globalenv prog_adc) m fd vargs t m' vres ->
    proc_state_related (of_mem proc m') e 
    (unpredictable Arm6_Message.EmptyMessage semstt).

(* Assume function reg_n only load from memory, not change it*)
Axiom get_reg_ok :
  forall e id m t m' r,
    eval_expr (Genv.globalenv prog_adc) e m RV (reg_id id) t m' r ->
    eval_expr (Genv.globalenv prog_adc) e m RV (reg_id id) t m r/\m=m'. 

Definition oldrn_assgnt := 
  Eassign (Evar old_Rn T1) (reg_id n) T1.

(* Assum the assignment of old_Rn has no effect on the part of memory
   where located proc*)
Axiom set_oldrn_ok:
  forall m m' v oldrn_blk ofs,
    store_value_of_type T1 m oldrn_blk ofs v = Some m'->
    of_mem proc m = of_mem proc m'.

Lemma oldrn_assgnt_ok:
 forall e m l b s t m' v,
  proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
  eval_expression (Genv.globalenv prog_adc) e m
    oldrn_assgnt t m' v ->
  proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)).
Proof.
  intros until v. intros psrel rn_as.
  inv rn_as. inv H. inv H4.
  eapply get_reg_ok in H5. inv H5.
  simpl in *.
  eapply set_oldrn_ok in H11.
  rewrite <- H11. exact psrel.
Qed.

(* Lemmas on if ConditionPassed*)
Definition condpass :=
  (Ecall (Evalof (Evar ConditionPassed T5) T5)
    (Econs
      (Eaddrof
        (Efield (Ederef (Evalof (Evar proc T3) T3) T6) cpsr
          T7) T8)
      (Econs (Evalof (Evar adc_compcert_fixed.cond T9) T9)
        Enil)) T4).

Axiom no_effect_condpass :
  forall e m m' t v,
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->    
    m = m'/\eval_expression (Genv.globalenv prog_adc) e m condpass t m' v.

Lemma condpass_false :
  forall m0 m0' e m t m' v cond s,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->
    Csem.is_false v T4 ->
    Arm6_Functions.State.ConditionPassed s cond = false.
Proof.
  intros until s. intros av cdps cdps_false.
  inv cdps_false.
  inv cdps. inv H. inv H0.
  inv H4. inv H3. inv H5. inv H3. inv H4. inv H14. inv H3. inv H4. inv H13.
  inv H3. inv H4. inv H10.
  inv H6.
  inv av. inv H14. inv H17. inv H18. inv H19. inv H20. inv H21. inv H22.
  pose (e:=
    (PTree.set old_Rn (b6, Tint I32 Unsigned)
      (PTree.set shifter_operand (b5, Tint I32 Unsigned)
        (PTree.set n (b4, Tint I8 Unsigned)
          (PTree.set d (b3, Tint I8 Unsigned)
            (PTree.set adc_compcert_fixed.cond 
              (b2, Tint I32 Signed)
              (PTree.set S (b0, Tint I8 Unsigned)
                (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                  empty_env)))))))).
  fold e in H7, H1.
  inv H1. unfold e in H6; simpl in H6; discriminate H6.
  inv H5. inv H10.
  (*to be improve *)
Qed.

Lemma condpass_true :
  forall m0 m0' e m t m' v cond s,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->
    Csem.is_true v T4 ->
    Arm6_Functions.State.ConditionPassed s cond = true.
Proof.
  intros until s. intros av cdps cdps_true.
  inv cdps. inv H. inv H4. inv H9. inv H5. inv H4. inv H5. inv H15. inv H4.
  inv H5. inv H14. inv H4. inv H5. inv H13.
  inv H0. inv H6.
  inv av. inv H14. inv H17. inv H18. inv H19. inv H20. inv H21. inv H22.
  pose (e:=
    (PTree.set old_Rn (b6, Tint I32 Unsigned)
      (PTree.set shifter_operand (b5, Tint I32 Unsigned)
        (PTree.set n (b4, Tint I8 Unsigned)
          (PTree.set d (b3, Tint I8 Unsigned)
            (PTree.set adc_compcert_fixed.cond 
              (b2, Tint I32 Signed)
                        (PTree.set S (b0, Tint I8 Unsigned)
                          (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                            empty_env)))))))).
  fold e in H7, H1.
  inv H1. unfold e in H6; simpl in H6; discriminate H6. inv H5. inv H10.
Qed.

(*Lemma on proc_state_relates holds after set_reg*)
Definition set_regpc :=
  Ecall (Evalof (Evar set_reg_or_pc T10) T10)
  (Econs (Evalof (Evar proc T3) T3)
    (Econs (Evalof (Evar d T4) T4)
      (Econs
        (Ebinop Oadd
          (Ebinop Oadd
            (Evalof (Evar old_Rn T1) T1)
            (Evalof (Evar shifter_operand T1) T1)
            T1)
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T4) T9)
          T9) Enil))) T11.

Lemma same_setregpc :
  forall e m l b s0 s t m' v d n so ,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    eval_expression (Genv.globalenv prog_adc) e m set_regpc t m' v ->
    (forall l b, proc_state_related (of_mem proc m') e 
      (Ok tt (mk_semstate l b
        (Arm6_State.set_reg s d (add (add (Arm6_State.reg_content s0 n) so)
          ((Arm6_State.cpsr s)[Cbit]) ))))).
Proof.
  intros until so. intros psrel setreg. intros.
  inv setreg. inv H. inv H4. inv H9. inv H5. inv H4. inv H5.
  inv H14. inv H4. inv H5. inv H13. inv H4. inv H17. inv H15. inv H4.
  inv H19. inv H4. inv H18. inv H4. inv H15. inv H13. inv H4. inv H5.
  inv H14. inv H0.
  (*inv H15.
  inv H4. inv H14. inv H19. inv H4. inv H18. inv H4. inv H14.
  inv H13. inv H4. inv H5.
  apply (functions_behavior_ok e l b s vf fd m2 vargs t3 m' vres l0 b0
    (Arm6_State.set_reg s d
      (add (add (Arm6_State.reg_content s0 n) so)
        (Arm6_State.cpsr s) [Cbit])))
    in psrel;
    [apply psrel|exact H11|exact H16].*)
Admitted.

(* Lemmas on if S==1 *)
Definition is_S_set :=
  Ebinop Oeq (Evalof (Evar S T4) T4)
  (Eval (Vint (repr 1)) T9) T9.

Lemma no_effect_is_S_set :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v ->
    m = m'/\eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v.
Proof.
  intros until v. intros is_s.
  split. inv is_s. inv H. inv H10. inv H4. inv H11. reflexivity. exact is_s.
Qed.

Lemma S_not_set:
  forall e m t m' v sbit,
    sbit_func_related m e sbit ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v ->
    Csem.is_false v T9 ->
    Util.zeq sbit 1 = false.
Proof.
  intros until sbit. intros sfrel s_set is_false. inv is_false.
  inv s_set. inv H. inv H10. inv H4. inv H11.
  inv H0. inv H7.
  inv sfrel.
  unfold bit_proj.
  unfold param_val. inv H5. inv H6. inv H2. rewrite H6.
  rewrite H7. unfold varg_proj.
  destruct v1; try auto.
    unfold sem_cmp in H0. unfold T4, T7, classify_cmp in H0. unfold typeconv in H0. 
    simpl in H0. unfold Val.of_bool in H0.
    unfold w1. 
    inv H0. destruct (eq i (repr 1)). inv H1. auto.
  rewrite H4. unfold varg_proj. simpl. reflexivity. 
Qed.

Lemma S_is_set:
  forall e m t m' v sbit,
    sbit_func_related m e sbit ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v ->
    Csem.is_true v T9 ->
    Util.zeq sbit 1 = true.
Proof.
  intros until sbit. intros sfrel s_set is_true.
  inv s_set. inv H. inv H10. inv H4. inv H11.
  inv H0. inv H6. inv H5. inv sfrel.
  simpl in H7.
  unfold bit_proj. unfold param_val. 
  inv H1.
    rewrite H6. rewrite H4. unfold varg_proj.
    destruct v1; 
      unfold sem_cmp in H7; unfold classify_cmp, T4, T7 in H7; simpl in H7; inv H7.
      inv is_true0. 
      assert (w1 = repr 1). auto. rewrite H0.
      unfold Val.of_bool in H. unfold Vtrue in H. unfold Vfalse in H.
      destruct (eq i (repr 1)). 
        inv H. simpl. reflexivity.
        inv H. induction H1. reflexivity.
      unfold Val.of_bool in H0.
      destruct (eq i (repr 1)). inv H0. inv H0.
    inv H5.
Qed.

(* Lemmas on if (((S == 1) && (d == 15)))*)
Definition is_S_set_and_is_pc :=
  Econdition
  (Ebinop Oeq (Evalof (Evar S T4) T4)
    (Eval (Vint (repr 1)) T9) T9)
  (Econdition
    (Ebinop Oeq (Evalof (Evar d T4) T4)
      (Eval (Vint (repr 15)) T9) T9)
    (Eval (Vint (repr 1)) T9)
    (Eval (Vint (repr 0)) T9) T9)
  (Eval (Vint (repr 0)) T9) T9.

Lemma no_effect_is_S_set_and_is_pc :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v ->
    m = m'/\eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v.
Proof.
  intros until v. intros spc. split.
  inv spc. inv H. inv H5. inv H13. inv H4. inv H16. inv H10.
  inv H4. inv H17. inv H4. inv H20. inv H12. reflexivity.
  inv H12. inv H4. inv H16. inv H4. inv H17. reflexivity.
  inv H10. inv H5. inv H12. inv H4. inv H13. reflexivity.
  exact spc.
Qed.

Lemma same_reg_val :
forall x y,
(eq x (repr y) = Util.zeq (mk_regnum x) y).
Proof.
Admitted.

Lemma S_set_and_is_pc_true:
  forall e m t m' v sbit d,
    sbit_func_related m e sbit ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v ->
    Csem.is_true v T9 ->
    Util.zeq sbit 1 && Util.zeq d 15 = true.
Proof.
  intros until d. intros sfrel dfrel spc spc_true.
  inv spc; inv H; simpl in *;
    (*true*)
    inv H5; inv H13; inv H4; inv H16; inv H6; inv H8.
    inv H7; inv H5; inv H3; simpl in H4.
      (*S exists*)
      inv sfrel; unfold bit_proj; unfold param_val. rewrite H8; rewrite H7.
      unfold varg_proj.
      destruct v2; simpl; try auto;
      unfold sem_cmp in H1; simpl in H1; inv H1.
      (*S is int*)
      unfold Val.of_bool in H9; unfold w1.
      destruct (eq i (repr 1)); simpl;
        [idtac|inv H9;destruct H2;reflexivity].
      (*S is set*)
      inv H10;
        (*d is 15*)
        simpl in H13; inv H16; inv H5; inv H18; inv H5;
        inv H19; inv H14; inv H20; inv H0; inv H6; inv H10; inv H5. 
        inv H1.
          (*d exists*)
          inv dfrel; unfold reg_proj; unfold param_val.
          rewrite H10. rewrite H6.
          unfold varg_proj.
          destruct v0;
          unfold sem_binary_operation in H11; simpl in H11;
          unfold sem_cmp in H11; simpl in H11; inv H11.
          (*d is int*)
          unfold Val.of_bool in H13.
          rewrite <- (same_reg_val i0).
          destruct (eq i0 (repr 15)). 
          reflexivity. inv H13; destruct H1; reflexivity.
          (*d not exist*)
          inv H5.
      (*S not set*)
      inv H1;
        (*d exists*)
        unfold sem_binary_operation in H11; unfold sem_cmp in H11; simpl in H11.
        inv dfrel; unfold reg_proj; unfold param_val.
        rewrite H10; rewrite H6.
        unfold varg_proj.
        destruct v0; inv H11. 
        (*d is int*)
          inv spc_true; destruct H1; auto.
        (*d not exist*)
        inv H5.
      (*S not exist*)
      inv H6.
    (*false*)
    inv H10; inv H0. inv H5. inv H7. inv H2.
      (*S exist*)
      inv sfrel; unfold bit_proj; unfold param_val. 
      rewrite H7; rewrite H6.
      unfold varg_proj.
      destruct v2; simpl; try auto;
      unfold sem_cmp in H1; simpl in H1; inv H1.
      (*i is int*)
      unfold Val.of_bool in H9; unfold w1.
      destruct (eq i (repr 1)); simpl.
        inv H9.
        inv H14. inv spc_true; destruct H1; auto.
      (*S not exist*)
      inv H5.  
Qed.        

Lemma S_set_and_is_pc_false:
  forall e m t m' v sbit d,
    sbit_func_related m e sbit ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v ->
    Csem.is_false v T9 ->
    Util.zeq sbit 1 && Util.zeq d 15 = false.
Proof.
  intros until d. intros sfrel dfrel spc spc_false.
  inv spc.
  inv H; simpl in *;
    (*true*)
    inv H5; inv H13; inv H4; inv H16; inv H6; inv H8.
    inv H7; inv H5; inv H3; simpl in H4.
      (*S exists*)
      inv sfrel; unfold bit_proj; unfold param_val; 
      rewrite H8; rewrite H7;
      unfold varg_proj.
      destruct v2; simpl; try auto;
      unfold sem_cmp in H1; simpl in H1; inv H1.
      (*v2 is int*)
      unfold Val.of_bool in H9; unfold w1.
      destruct (eq i (repr 1)); simpl;
        [idtac|inv H9;destruct H2;reflexivity].
        (*i is false*)
        inv H10;
        simpl in H13; inv H16; inv H5; inv H18; inv H5;
        inv H19; inv H14; inv H20; inv H0; inv H6; inv H10; inv H5. 
        (*d is 15*)
        inv spc_false.
        (*d is not 15*)
        inv H1.
          (*d exists*)
          unfold sem_binary_operation in H11; simpl in H11;
          unfold sem_cmp in H11; simpl in H11; inv H11.
          inv dfrel; unfold reg_proj; unfold param_val; unfold varg_proj.
          rewrite H10; rewrite H6.
          destruct v0; inv H0.
            (*d is int*)
            unfold Val.of_bool in H13.
            rewrite <- (same_reg_val i0).
            destruct (eq i0 (repr 15)). inv H13. reflexivity.
          (*d not exist*)
          inv H5.
      (*S not exist*)
      inv H6.
    (*false*)
    inv H10. inv H0. inv H14. inv H7. inv H5.
    inv H2.
      (*S exists*)
      inv sfrel; unfold bit_proj; unfold param_val; unfold varg_proj.
      rewrite H7; rewrite H6.
      destruct v2; inv H1.
      (*S is int*)
      unfold Val.of_bool in H9. unfold w1.
      destruct (eq i (repr 1)). inv H9. auto.
      (*S not exist*)
      inv H5.
Qed.

(* Lemmas on if CurrentModeHasSPSR *)
Definition hasSPSR :=
  Ecall (Evalof (Evar CurrentModeHasSPSR T12) T12)
  (Econs (Evalof (Evar proc T3) T3) Enil) T4.

Axiom if_hasSPSR_ok :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    m = m'/\eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v.

Lemma hasSPSR_true' :
  forall m0 m0' e m vargs t m' v l b s,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)) ->
    Csem.is_true v T4 ->
    word_of_proc_mode (mode_proj m' e) < 5.
Proof.
  intros until s. intros av bp hs psrel tr.

  inv hs. inv H. inv H0. 
  (* m = m3 *)
  inv H4. inv H3. inv H5. inv H3. inv H4. inv H13.
  (* ? *)
  inv H6.
  (* expand local env e *)
  inv av. inv H14. inv H17. inv H18. inv H19. inv H20. inv H21. inv H22.
  pose (e:=
    PTree.set old_Rn (b7, Tint I32 Unsigned)
      (PTree.set shifter_operand (b6, Tint I32 Unsigned)
        (PTree.set n (b5, Tint I8 Unsigned)
          (PTree.set d (b4, Tint I8 Unsigned)
            (PTree.set cond (b3, Tint I32 Signed)
              (PTree.set S (b2, Tint I8 Unsigned)
                (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                  empty_env))))))).
  fold e in psrel, bp, H7. fold e. 
  (* CurrentModeHasSPSR is in global env *)
  inv H1; [simpl in H6; discriminate H6| clear H3].
  (* search CurrentModeHasSPSR in global env *)
  (* vf=Vptr (-6) w0 *)
  inv H5. unfold load_value_of_type in H4; simpl in H4. 
  injection H4; intro; clear H4. rewrite <- H in *; clear vf H.
  (* fd = fun_Internal_CurrentModeHasSPSR *)
  inversion H11;  destruct eq_dec; 
    [clear e0 H11 H2 H12 H8; inv H0|discriminate H0].

  (* pass parameter proc to internal function CurrentModeHasSPSR *)
  inv H7. inv H5. 
  (* v0 is value of proc *)
  inv H1; clear H4.
  inv H3;
  [unfold e in H5;simpl in H5;injection H5;intro;rewrite<-H in *;clear b0 H H5
  |unfold e in H1;simpl in H1;discriminate H1].


  (* open CrrentModeHasSPSR *)
  inv H16. inv H4. 
  (* return value is v (cast from v1) *)
  simpl in H5; destruct H5.
  (* m9 = m10 *)
  inv H11. inv H5. inv H27. inv H26. inv H16. inv H25. inv H24. inv H16. inv H21.
  (* arguments v2,v3 of binary operation lt*)
  inv H7. simpl in H23.
  (* v3 = 5 *)
  inv H22.
  (* v2 = v0 *)
  inv H21; clear H11.
  (* typ_struct_SLv6_StatusRegister is a structure *)
  inv H9;[idtac|simpl in H24;unfold T7 in H24;discriminate H24].
  inv H24.
  (* offset of mode is 16 *)
  assert (field_offset mode typ_struct_SLv6_StatusRegister = OK 16).  
  unfold field_offset. simpl. 
  Ltac unfold_identeq :=
    destruct AST.ident_eq;
      [try (unfold align;simpl;discriminate||destruct AST.ident_eq)
        |try unfold_identeq].
  unfold_identeq. unfold align. simpl. reflexivity. admit.
  rewrite H5 in H25; clear H5. 
  injection H25;intro;rewrite<-H5 in H16;clear H5 H25 delta.
  (* typ_struct_SLv6_Processor is a structure *)    
  inv H12; [idtac|simpl in H24;unfold T6 in H24;discriminate H24].
  inv H24.
  (* offset of cpsr  is 2 *)
  assert (field_offset cpsr typ_struct_SLv6_Processor = OK 2). admit.
  rewrite H5 in H25; clear H5. 
  injection H25; intro; rewrite<-H5 in H16; clear delta H5 H25.
  (* expand e0 *)
  inv H1. inv H26.   
  (* proc is in e0 *)
  inv H11. inv H12. inv H7;[idtac|simpl in H11; discriminate H11]. clear H9.
  (* b9 = b8 *)
  simpl in H22; injection H22;intro;rewrite<-H1 in *; clear b9 H22 H1.
  (* load v0 from b9 *)
  inv H3.
  inv H28; simpl in H26;injection H26;intro;rewrite<-H1 in *;clear b9 H1 H26.
  unfold store_value_of_type in H27;simpl in H27.
  generalize H27; intro bp'.
  apply Mem.load_store_same in H27;
    [idtac|simpl;destruct v0;simpl;try(exact I||inv H2)].
  unfold load_value_of_type in *; simpl in H6, H16, H21.
  rewrite H27 in H21. 
  injection H21; intro. destruct v0; try discriminate H1.
  injection H1; intros; rewrite<-H3,H5 in *;clear H1 H3 H5.
  simpl in H27.
  (* v' = Vptr b0 i*)
  inv H2.
  unfold sem_cmp in H23; simpl in H23.
  destruct v2; try discriminate H23.
  injection H23; intro; clear H23. rewrite <- H1 in *; clear H1.

  (* unfold goal *)
  unfold mode_proj. unfold find_mode. unfold find_cpsr. unfold find_field.
  unfold proc_loc. 
  unfold e. Set Printing Depth 50. simpl. unfold load_value_of_type; simpl.
  (* b1 not change between m3 m8 *)
  generalize H6;intro.
  apply (Mem.load_alloc_other m3 0 (sizeof (Tpointer typ_SLv6_Processor))
    m8 b8 H25) in H6. 
  (* b1 not changed between m8 m10 *)
  (*apply load_store*)
Admitted.

Lemma hasSPSR_true :
  forall m0 m0' m0'' e m vargs t m' v l b s em,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m0'' ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)) ->
    Csem.is_true v T4 ->
    Arm6_State.mode s = exn  em.
Proof.
  intros until em. intros av bp hs psrel tr.
  inv hs. inv H. inv H0. inv H4. inv H3. inv H5. inv H3. inv H4. inv H13.
  inv H6.
  inv av. inv H14. inv H17. inv H18. inv H19. inv H20. inv H21. inv H22.
  pose (e:=
    PTree.set old_Rn (b7, Tint I32 Unsigned)
            (PTree.set shifter_operand (b6, Tint I32 Unsigned)
               (PTree.set n (b5, Tint I8 Unsigned)
                  (PTree.set d (b4, Tint I8 Unsigned)
                     (PTree.set cond (b3, Tint I32 Signed)
                        (PTree.set S (b2, Tint I8 Unsigned)
                           (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                              empty_env))))))).
  fold e in psrel, bp, H7. inv H1. simpl in H6; discriminate H6. simpl in H3.
  inv H5. inv H4. inv H11. 
  destruct eq_dec; [clear e0|discriminate H0].
  clear H2 H12. inv H0. inv H7. inversion H8; clear H8. 
  rewrite <- H0 in *; clear H0. rewrite <- H4 in *; clear H4. clear H5.
  inv H6.
  
  inv H1. clear H5. 
  inv H4; [idtac|unfold e in H1; simpl in H1; discriminate H1].
  unfold e in H6; simpl in H6; inversion H6. rewrite <- H0 in *; clear b0 H0 H6.
  unfold load_value_of_type in H7; simpl in H7.

  (* open CrrentModeHasSPSR *)
  inv H16. inv H5. simpl in H6. destruct H6.

Admitted.

Lemma hasSPSR_false :
  forall e m t m' v s,
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    Csem.is_false v T4 ->
    Arm6_State.mode s = usr.
Proof.
Admitted.

(*Lemma on proc_state_relates holds after copy_StatusRegister*)
Definition get_spsr :=
  Ecall (Evalof (Evar spsr T14) T14)
  (Econs (Evalof (Evar proc T3) T3)
    Enil) T8.

Axiom get_spsr_ok:
  forall e m t m' r,
    eval_expr (Genv.globalenv prog_adc) e m RV get_spsr t m' r ->
    m = m'.

Definition cp_SR :=
  Ecall
  (Evalof (Evar copy_StatusRegister T13) T13)
  (Econs
    (Eaddrof
      (Efield
        (Ederef (Evalof (Evar proc T3) T3) T6)
        cpsr T7) T8)
    (Econs
      (Ecall (Evalof (Evar spsr T14) T14)
        (Econs (Evalof (Evar proc T3) T3)
          Enil) T8) Enil)) T11.

Lemma same_cp_SR :
  forall e m l b s t m' v em,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    eval_expression (Genv.globalenv prog_adc) e m cp_SR t m' v ->
    (forall l b, proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b
      (Arm6_State.set_cpsr s (Arm6_State.spsr s em))))).
Proof.
  intros until em. intros psrel cpsr l' b'.
  inv cpsr. inv H. inv H4. inv H9. simpl in *.
  inv H5. inv H4. inv H5. inv H15. inv H4. inv H5.
  inv H14. inv H4. inv H3. inv H15. inv H5. inv H4. inv H5. inv H21.
  inv H13. simpl in *.
  (* Function spsr, get spsr from the current state *)
  apply (functions_behavior_ok e l b s vf0 fd0 m4 vargs0 t5 m2 vres0 l b s) 
    in psrel; [idtac|exact H18|exact H23].
  (* Function copy_StatusRegister, copy the current spsr to cpsr*)
  apply (functions_behavior_ok e l b s vf fd m2 vargs t3 m' vres l' b'
    (Arm6_State.set_cpsr s (Arm6_State.spsr s em)))
    in psrel; [idtac|exact H11|exact H16].
  exact psrel.
Qed.

(* Lemma on proc_state_relates holds after unpredictable*)
(* In fact, unpredictable in simlight is a annotation, which will print
   a error message. 
   For the moment, we consider it as a function call with an 
   empty body *)
Definition unpred :=
  (Ecall (Evalof (Evar unpredictable T15) T15) Enil T11).

Lemma same_unpred :
  forall e m s t m' v,
    proc_state_related (of_mem proc m) e (Ok tt s) ->
    eval_expression (Genv.globalenv prog_adc) e m unpred t m' v ->
    proc_state_related (of_mem proc m') e (Ko Arm6_Message.EmptyMessage).
Proof.
  intros until v. intros psrel unp.
  inv unp. inv H. inv H4. inv H9. inv H5.
  apply (funct_unpredictable e s vf fd m2 vargs t3 m' vres) in psrel;
  unfold unpredictable in psrel; unfold raise in psrel; 
  [exact psrel|exact H11|exact H16].
Qed.

(* Lemma on proc_state_relates holds after NZCV flag setting*)
Definition nflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef (Evalof (Evar proc T3) T3) T6)
      cpsr T7) N_flag T4)
  (Ecall (Evalof (Evar get_bit T16) T16)
    (Econs
      (Ecall (Evalof (Evar reg T2) T2)
        (Econs (Evalof (Evar proc T3) T3)
          (Econs 
            (Evalof (Evar d T4) T4) Enil))
        T1)
      (Econs (Eval (Vint (repr 31)) T9)
        Enil)) T4) T4.

Lemma same_nflag_assgnt :
  forall e m l b s d t m' v,
  proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
  d_func_related m e d ->
  eval_expression (Genv.globalenv prog_adc) e m nflag_assgnt t m' v->
  forall l b,
  proc_state_related (of_mem proc m') e
    (Ok tt
        (mk_semstate l b
           (Arm6_State.set_cpsr_bit s Nbit
              (Arm6_State.reg_content s d) [n31] )
         )
    ).
Proof.
Admitted.

Definition zflag_assgnt :=
  Eassign
  (Efield
    (Efield
      (Ederef 
        (Evalof (Evar proc T3) T3) T6)
      cpsr T7) Z_flag T4)
  (Econdition
    (Ebinop Oeq
      (Ecall (Evalof (Evar reg T2) T2)
        (Econs
          (Evalof (Evar proc T3) T3)
          (Econs
            (Evalof (Evar d T4) T4)
            Enil)) T1)
      (Eval (Vint (repr 0)) T9) T9)
    (Eval (Vint (repr 1)) T9)
    (Eval (Vint (repr 0)) T9) T9) T4.

Lemma same_zflag_assgnt :
  forall e m l b s d t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m zflag_assgnt t m' v->
    forall l b, proc_state_related (of_mem proc m') e 
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Zbit
        (if Util.zeq (Arm6_State.reg_content s d) 0
         then repr 1
         else repr 0)))).
Proof.
Admitted.

Definition cflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef
        (Evalof (Evar proc T3) T3)
        T6) cpsr T7) C_flag T4)
  (Ecall
    (Evalof 
      (Evar CarryFrom_add3 T17) T17)
    (Econs
      (Evalof (Evar old_Rn T1) T1)
      (Econs
        (Evalof
          (Evar shifter_operand T1)
          T1)
        (Econs
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T4) T4)
          Enil))) T4) T4.

Lemma same_cflag_assgnt:
  forall m e l b s0 s n so t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    n_func_related m e n ->
    so_func_related m e so ->
    eval_expression (Genv.globalenv prog_adc) e m cflag_assgnt t m' v->
    forall l b, proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Cbit
        (Arm6_Functions.CarryFrom_add3 (Arm6_State.reg_content s0 n) so
          (Arm6_State.cpsr (st (mk_semstate l b s))) [Cbit])))).
Proof.
Admitted.

Definition vflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef
        (Evalof (Evar proc T3) T3)
        T6) cpsr T7) V_flag T4)
  (Ecall
    (Evalof
      (Evar OverflowFrom_add3 T18)
      T18)
    (Econs
      (Evalof (Evar old_Rn T1) T1)
      (Econs
        (Evalof
          (Evar shifter_operand T1)
          T1)
        (Econs
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T4) T4)
          Enil))) T4) T4.

Lemma same_vflag_assgnt:
  forall m e l b s0 s n so t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    n_func_related m e n ->
    so_func_related m e so ->
    eval_expression (Genv.globalenv prog_adc) e m vflag_assgnt t m' v->
    proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Arm6_SCC.Vbit
        (Arm6_Functions.OverflowFrom_add3 (Arm6_State.reg_content s0 n) so
           (Arm6_State.cpsr (st (mk_semstate l b s))) [Cbit])))).
Proof.
Admitted.


(* During function execution, none other parameters are changed*)
Lemma cp_SR_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m cp_SR Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma reg_S_not_changed :
  forall e m vargs t m' v,
    eval_funcall (Genv.globalenv prog_adc) m (Internal fun_internal_reg) 
    vargs t m' v ->
    param_val S m e = param_val S m' e.
Proof.
Admitted.


Lemma diff_block :
  forall m1 ofs1 b1 m2 ofs2 b2 m3,
    Mem.alloc m1 0 ofs1 = (m2, b1) ->
    Mem.alloc m2 0 ofs2 = (m3, b2) ->
    b1 < b2.
Proof.
  intros until m3. intros alc1 alc2.
  apply Mem.valid_new_block in alc1. unfold Mem.valid_block in alc1.
  apply Mem.alloc_result in alc2. rewrite <- alc2 in alc1. exact alc1.
Qed.


Lemma rn_ass_S_not_changed:
  forall m0 m0' vargs m e v m', 
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    list_norepet 
    (var_names fun_internal_ADC.(fn_params) ++ var_names fun_internal_ADC.(fn_vars)) ->
    eval_expression (Genv.globalenv prog_adc) e m oldrn_assgnt Events.E0 m' v ->
    param_val S m e = param_val S m' e.
Proof.
  intros until m'. intros av bp ln evex.
  unfold param_val.
  inv bp. inv H8. rewrite H5.
  inv H11. inv H13. inv H15. inv H17. inv H19.
  unfold store_value_of_type in *. simpl in H7, H10, H12, H14, H16, H18.

  inv av. 
  inv H19. inv H21. inv H22. inv H23. inv H24. inv H25. inv H26.
  simpl in H4, H5, H6, H8, H9, H11.
  inv H4. inv H5. inv H6. inv H8. inv H9. inv H11. 

  assert (lt01:b0 < b1).
  apply (diff_block m7 (sizeof (Tint I8 Unsigned)) b0) in H19;
    [exact H19| exact H20].

  assert (lt12:b1 < b2).
  apply (diff_block m8 (sizeof (Tint I32 Signed)) b1) in H21;
    [exact H21| exact H19].

  assert (lt23:b2 < b3).
  apply (diff_block m9 (sizeof (Tint I8 Unsigned)) b2) in H22;
    [exact H22| exact H21].

  assert (lt34:b3 < b4).
  apply (diff_block m10 (sizeof (Tint I8 Unsigned)) b3) in H23;
    [exact H23| exact H22].

  assert (lt411:b4 < b11).
  apply (diff_block m11 (sizeof (Tint I32 Unsigned)) b4) in H24;
    [exact H24| exact H23].

  generalize lt34; intro.
  apply (Zlt_trans b2) in lt0;
    [apply (Zlt_trans b1) in lt0; 
      [apply (Zlt_trans b0) in lt0;[idtac|exact lt01] |exact lt12]|exact lt23].
  
  assert (load_value_of_type (Tint I8 Unsigned) m4 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m3 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m3 b1 (signed w0) v2);
    [exact H12 | left; apply Zlt_not_eq in lt01; exact lt01].
    
  assert (load_value_of_type (Tint I8 Unsigned) m5 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m4 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint8unsigned m4 b2 (signed w0) v3);
    [exact H14|left; apply (Zlt_trans b0) in lt12;
                       [apply Zlt_not_eq in lt12;exact lt12|exact lt01]].

  assert (load_value_of_type (Tint I8 Unsigned) m6 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m5 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint8unsigned m5 b3 (signed w0) v4);
    [exact H16|left; apply (Zlt_trans b1) in lt23;
                       [apply (Zlt_trans b0) in lt23;
                         [apply Zlt_not_eq in lt23;
                           exact lt23|exact lt01]|exact lt12]].

  assert (load_value_of_type (Tint I8 Unsigned) m b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m6 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m6 b4 (signed w0) v5);
    [exact H18|left;apply (Zlt_trans b2) in lt34;
                      [apply (Zlt_trans b1) in lt34;
                         [apply (Zlt_trans b0) in lt34;
                            [apply Zlt_not_eq in lt34;
                              exact lt34|exact lt01]|exact lt12]|exact lt23]].

  rewrite <- H2 in H1; clear H2.
  rewrite <- H1 in H0; clear H1.
  rewrite <- H0 in H; clear H0.
  
  rename H24 into alc12, H17 into alc0, H20 into alc7, H19 into alc8, H21 into alc9,
    H22 into alc10, H23 into alc11.
  rename H7 into st0, H10 into st2, H12 into st3, H14 into st4, H16 into st5,
    H18 into st6.
  rename H into Heqmm3.
  pose (e:=(PTree.set old_Rn (b11, Tint I32 Unsigned)
              (PTree.set shifter_operand (b4, Tint I32 Unsigned)
                 (PTree.set n (b3, Tint I8 Unsigned)
                    (PTree.set d (b2, Tint I8 Unsigned)
                       (PTree.set cond (b1, Tint I32 Signed)
                          (PTree.set S (b0, Tint I8 Unsigned)
                             (PTree.set proc (b, Tpointer typ_SLv6_Processor)
                                empty_env)))))))).
  fold e in evex.
  
  (* begin with assgn expr *)
  inv evex. inv H. inv H0.
  inv H5. inv H6. inv H10. inv H2. inv H10.
  inv H3. inv H6. inv H3. inv H18. inv H3. inv H6. inv H14.
  clear H15 H9.

  (* reg is in loc env *)
  assert (reg_not_loc: e!reg = None).
  unfold e. simpl. reflexivity.
  inv H5. inv H1. rewrite reg_not_loc in H9. discriminate H9. clear H3.

  (* ofs is w0 *)
  inv H5. clear H2. inv H6. inv H16.
  destruct eq_dec; [idtac|discriminate H0]. clear e0. inv H0.

  (*
  (* open internal function reg *)
  inv H21. inv H1. inv H20. inv H21.

  (* nextblock is not change from Mem.store on memory *)
  generalize alc12; intro.
  apply Mem.valid_new_block in alc1. unfold Mem.valid_block in alc1.
  apply Mem.nextblock_store in st0.
  apply Mem.nextblock_store in st2.
  apply Mem.nextblock_store in st3.
  apply Mem.nextblock_store in st4.
  apply Mem.nextblock_store in st5.
  apply Mem.nextblock_store in st6.
  rewrite <- st6 in st5. rewrite <- st5 in st4. rewrite <- st4 in st3. 
  rewrite <- st3 in st2. rewrite <- st2 in st0.
  rewrite <- st0 in alc1.

  (* b0 < b6 *)
  generalize H19; intros.
  apply Mem.alloc_result in H19. rewrite <- H19 in alc1.
  apply (Zlt_trans b4) in alc1; [idtac|exact lt411]. 
  apply (Zlt_trans b0) in alc1; [idtac|exact lt0].

  (* expand bind_parameters *)
  inv H2. inv H23. inv H24. simpl in H16, H15.
  inversion H16. rewrite <- H2 in *. clear b8 H16 H2.
  inversion H15. rewrite H2 in *. clear b7 H15 H2.

  (* between m15 and m17 *)  
  assert (load_value_of_type (Tint I8 Unsigned) m17 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m15 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_alloc_unchanged m15 0 
    (sizeof (Tpointer typ_SLv6_Processor)) m17 (Mem.nextblock m15));
  [exact H1|unfold Mem.valid_block; exact alc1].
  
  (* between m17 and m1 *)
  generalize H18; intro.
  apply Mem.valid_new_block in H1. unfold Mem.valid_block in H1.
  apply Mem.alloc_result in H18.
  apply (Zlt_trans b0) in H1; [idtac|exact alc1].
  assert (load_value_of_type (Tint I8 Unsigned) m1 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m17 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_alloc_unchanged m17 0 
    (sizeof (Tint I8 Unsigned)) m1 b6);
  [exact H2|unfold Mem.valid_block; exact H1].
  rewrite <- H6 in H. clear H6.

  (* between m1 and m18 *)
  unfold store_value_of_type in H22, H21; simpl in H22, H21.
  assert (load_value_of_type (Tint I8 Unsigned) m18 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m1 b0 w0). 
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m1 ((Mem.nextblock m15)) (signed w0) v7);
    [exact H22|left;apply Zlt_not_eq in alc1; exact alc1].
  rewrite <- H6 in H. clear H6.

  (* betwwen m18 and m13 *)
  assert (load_value_of_type (Tint I8 Unsigned) m13 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m18 b0 w0). 
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint8unsigned m18 b6 (signed w0) v8);
    [exact H21|left; apply Zlt_not_eq in H1; rewrite <- H18 in H1; exact H1].
  rewrite <- H6 in H. clear H6.

  (* between m13 and m16 *)
  pose (e0 := (PTree.set adc_compcert_fixed.reg_id (b6, Tint I8 Unsigned)
            (PTree.set proc (Mem.nextblock m15, Tpointer typ_SLv6_Processor)
               empty_env))).
  (*fold e0 in H3.
  inv H3. inv H15.*)
  inv H3. fold e0 in H15. inv H15.  inv H3. inv H16.
*)

  apply (reg_S_not_changed e m15 vargs t3 m14 v6) in H21.
  unfold param_val in H21. unfold e in H21; simpl in H21.
  unfold store_value_of_type in H12; simpl in H12.

  assert (Heqm'm14: load_value_of_type (Tint I8 Unsigned) m' b0 w0=
  load_value_of_type (Tint I8 Unsigned) m14 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m14 b5 (signed ofs) v). exact H12.
  left.
  inv H7; [idtac|inv H2]. 
  unfold e in H3; simpl in H3. inversion H3. rewrite <- H0 in *.
  clear b5 H0.
  apply (diff_block m11 (sizeof (Tint I32 Unsigned)) b4) in alc12;
    [apply (Zlt_trans b0) in alc12; 
      [apply Zlt_not_eq in alc12; exact alc12|exact lt0] |exact alc11].
  
  rewrite H21. rewrite Heqm'm14. reflexivity.
Qed.

Lemma rn_ass_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m oldrn_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma set_reg_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m set_regpc Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma unpred_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m unpred Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma nf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m nflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma zf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m zflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma vf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m vflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma cf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m cflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma same_bool : forall b, b&&b = b.
Proof.
  destruct b;simpl;reflexivity.
Qed.

Theorem related_aft_ADC: forall e m0 m1 m2 mfin vargs s out sbit cond d n so,
  alloc_variables empty_env m0 (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m1 ->
  bind_parameters e m1 fun_internal_ADC.(fn_params) vargs m2 ->
(* TODO: valid_access needs to be more precise *)
  (forall m ch b ofs, Mem.valid_access m ch b ofs Readable) ->
  proc_state_related (of_mem proc m2) e (Ok tt (mk_semstate nil true s)) ->
  sbit_func_related m2 e sbit ->
  cond_func_related m2 e cond ->
  d_func_related m2 e d ->
  n_func_related m2 e n ->
  so_func_related m2 e so ->
(* Comparison between eval_funcall, exec_stmt:
   [eval_funcall] is big step semantic. It can be seen as 6 steps, 
   and we can observe 4 times of memory changes.
   1. Check there are no repetitive parameters in function parameter list;
   2. Allocate function parameters into memory and fill them in the empty local environment (m0->m1);
   3. Bind these parameters with there initial values (m1->m2);
   4. Execute all the statement of the function body (m2->m3);
   5. Clean up the memory which are used to store the local parameters when
   execution finishes (m3->m4).
   This final memory doesn't contain the final [proc] we expect. It is in [m3], but in [m4],
   their memory blocks are freed.
   [exec_stmt] is also big step semantic. It indicates the outcome of 
   statement execution [Out_break], [Out_continue], [Out_normal] and [Out_return].
   The final memory state is the memory which contains the final values of parameters.
   The final [proc] is in this memory state which we want to relate.*)
  exec_stmt (Genv.globalenv prog_adc) e m2 fun_internal_ADC.(fn_body) Events.E0 mfin out ->
  proc_state_related (of_mem proc mfin) e (S.ADC_step sbit cond d n so (mk_semstate nil true s)). 
Proof.
  
  intros until so.
  intros al bi valacc psrel sfrel cfrel dfrel nfrel sofrel exstmt.

  inv exstmt; [idtac | nod];
  apply Events.Eapp_E0_inv in H3; destruct H3; subst.
  rename H4 into rn_assgnt, H7 into main_p.
  inv rn_assgnt;
  rename H2 into rn_assgnt.
  apply (oldrn_assgnt_ok e m2 nil true s Events.E0 m3 v) in psrel; 
    [idtac|exact rn_assgnt];
  unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 S) in sfrel;
    [idtac | exact rn_assgnt];
  fold (bit_proj m3 e S) in sfrel; fold (sbit_func_related m3 e sbit) in sfrel.
  unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert_fixed.cond) in cfrel;
    [idtac | exact rn_assgnt];
  fold (cond_proj m3 e) in cfrel; fold (cond_func_related m3 e cond) in cfrel.
  unfold d_func_related in dfrel; unfold reg_proj in dfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert_fixed.d) in dfrel;
    [idtac | exact rn_assgnt];
  fold (reg_proj m3 e adc_compcert_fixed.d) in dfrel; fold (d_func_related m3 e d) in dfrel.
  unfold n_func_related in nfrel; unfold reg_proj in nfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert_fixed.n) in nfrel;
    [idtac | exact rn_assgnt]; 
  fold (reg_proj m3 e adc_compcert_fixed.n) in nfrel; fold (n_func_related m3 e n) in nfrel.
  unfold so_func_related in sofrel; unfold bits_proj in sofrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 shifter_operand) in sofrel;
    [clear rn_assgnt | exact rn_assgnt];
  fold (bits_proj m3 e shifter_operand) in sofrel; fold (so_func_related m3 e so) in sofrel (* m2=m3 *).
  inv main_p;
  rename H5 into condpass, H8 into cp_b, H9 into main_p, H4 into evs;
      simpl in cp_b;
      apply Events.Eapp_E0_inv in evs; destruct evs; subst;
      apply no_effect_condpass in condpass0; 
      inversion condpass0 (* m3=m4 *);
      rewrite H in * |- *; clear H condpass0;
      rename H0 into condpass.
    (* ConditionPassed(&proc->cpsr, cond) evaluates to true *)
    apply (condpass_true m0 m1 e m4 Events.E0 m4 v1 cond s) in cp_b;
    [idtac| exact al| exact condpass].
      (*[idtac |exact al | inv cp_b].*)

    inv main_p; [idtac | nod];
    rename H4 into setreg, H7 into main_p, H3 into evs;
    apply Events.Eapp_E0_inv in evs; destruct evs; subst.

    inv setreg;
    rename H2 into setreg;
    apply (same_setregpc e m4 nil true s s Events.E0 m5 v0 d n so) 
      with nil (Util.zne d 15) in psrel;
      [idtac | fold set_regpc in setreg; apply setreg].
    unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
    rewrite (set_reg_params_not_changed m4 e v0 m5 S) in sfrel;
      [idtac | exact setreg];
    fold (bit_proj m5 e S) in sfrel; fold (sbit_func_related m5 e sbit) in sfrel.
    unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
    rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert_fixed.cond) in cfrel;
      [idtac | exact setreg];
    fold (cond_proj m5 e) in cfrel; fold (cond_func_related m5 e cond) in cfrel.
    unfold d_func_related in dfrel; unfold reg_proj in dfrel;
    rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert_fixed.d) in dfrel;
      [idtac | exact setreg];
    fold (reg_proj m5 e adc_compcert_fixed.d) in dfrel; fold (d_func_related m5 e d) in dfrel.
    unfold n_func_related in nfrel; unfold reg_proj in nfrel;
    rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert_fixed.n) in nfrel;
      [idtac | exact setreg]; 
    fold (reg_proj m5 e adc_compcert_fixed.n) in nfrel; fold (n_func_related m5 e n) in nfrel.
    unfold so_func_related in sofrel; unfold bits_proj in sofrel;
    rewrite (set_reg_params_not_changed m4 e v0 m5 shifter_operand) in sofrel;
      [clear setreg | exact setreg];
    fold (bits_proj m5 e shifter_operand) in sofrel; fold (so_func_related m5 e so) in sofrel (*m4 -> m5*).
    inv main_p;
    rename H5 into sd, H8 into sd_b, H9 into main_p, H4 into evs;
        simpl in sd_b;
        apply no_effect_is_S_set_and_is_pc in sd; 
        inversion sd; 
        rewrite H in * |- *; clear H sd; (* m5=m6 *)
        rename H0 into sd;
        apply Events.Eapp_E0_inv in evs; destruct evs; subst.
      (* ((S == 1) && (d == 15)) evaluates to true *)
      apply (S_set_and_is_pc_true e m6 Events.E0 m6 v2 sbit d) in sd;
        [idtac|exact sfrel|exact dfrel|exact sd_b].
      inv main_p;
      rename H5 into hasspsr, H8 into spsr_b, H9 into main_p, H4 into evs;
          simpl in spsr_b;
          apply Events.Eapp_E0_inv in evs; destruct evs; subst;
          apply if_hasSPSR_ok in hasspsr;
          inversion hasspsr;
          rewrite H in * |- *; 
          clear H hasspsr; rename H0 into hasspsr (* m6=m7*).
        (* CurrentModeHasSPSR(proc) evaluates to true *)
        inv main_p;
        rename H2 into cp_sr.
        generalize psrel; intro psrelm7.
        apply (same_cp_SR e m7 nil (Util.zne d 15) 
          (Arm6_State.set_reg s d
          (add (add (Arm6_State.reg_content s n) so)
            (Arm6_State.cpsr s) [Cbit])) Events.E0 mfin v4 und) 
        with nil (Util.zne d 15) in psrel;
          [idtac | exact cp_sr ].
        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (cp_SR_params_not_changed m7 e v4 mfin S) in sfrel;
          [idtac | exact cp_sr];
        fold (bit_proj mfin e S) in sfrel; fold (sbit_func_related mfin e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert_fixed.cond) in cfrel;
          [idtac | exact cp_sr];
        fold (cond_proj mfin e) in cfrel; fold (cond_func_related mfin e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert_fixed.d) in dfrel;
          [idtac | exact cp_sr];
        fold (reg_proj mfin e adc_compcert_fixed.d) in dfrel; fold (d_func_related mfin e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert_fixed.n) in nfrel;
          [idtac | exact cp_sr]; 
        fold (reg_proj mfin e adc_compcert_fixed.n) in nfrel; fold (n_func_related mfin e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (cp_SR_params_not_changed m7 e v4 mfin shifter_operand) in sofrel;
          [clear cp_sr | exact cp_sr];
        fold (bits_proj mfin e shifter_operand) in sofrel; fold (so_func_related mfin e so) in sofrel (*m7->mfin*).
        apply (hasSPSR_true m0 m1 m2 e m7 vargs Events.E0 m7 v3 nil (Util.zne d 15)
          (Arm6_State.set_reg s d
            (add (add (Arm6_State.reg_content s n) so)
              (Arm6_State.cpsr s) [Cbit]))
          und) in spsr_b;
          [idtac |exact al|exact bi|exact hasspsr|exact psrelm7].
        unfold S.ADC_step; unfold _get_st; unfold bind_s;
          unfold bind; simpl.
        rewrite cp_b; rewrite sd; simpl.
        unfold if_CurrentModeHasSPSR; unfold block; unfold fold_left;
        unfold _get_bo; unfold bind_s; unfold next; unfold bind; simpl;
        unfold _Arm_State.set_reg.
        rewrite spsr_b; simpl; unfold _Arm_State.set_reg; unfold _Arm_State.set_cpsr.
        unfold _set_bo; unfold ok_semstate. unfold loc. unfold st. rewrite same_bool.
        exact psrel. (*exact hasspsr. exact hasspsr.*)
        (* CurrentModeHasSPSR(proc) evaluates to false *)
        inv main_p; rename H2 into unp.
        apply (same_unpred e m7 
                (mk_semstate nil (Util.zne d 15) (Arm6_State.set_reg s d
                  (add (add (Arm6_State.reg_content s n) so)
                    (Arm6_State.cpsr s) [Cbit])))
                Events.E0 mfin v4) in psrel;
        [idtac | exact unp].
        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (unpred_params_not_changed m7 e v4 mfin S) in sfrel;
          [idtac | exact unp];
        fold (bit_proj mfin e S) in sfrel; fold (sbit_func_related mfin e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert_fixed.cond) in cfrel;
          [idtac | exact unp];
        fold (cond_proj mfin e) in cfrel; fold (cond_func_related mfin e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert_fixed.d) in dfrel;
          [idtac | exact unp];
        fold (reg_proj mfin e adc_compcert_fixed.d) in dfrel; fold (d_func_related mfin e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert_fixed.n) in nfrel;
          [idtac | exact unp]; 
        fold (reg_proj mfin e adc_compcert_fixed.n) in nfrel; fold (n_func_related mfin e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (unpred_params_not_changed m7 e v4 mfin shifter_operand) in sofrel;
          [clear unp | exact unp];
        fold (bits_proj mfin e shifter_operand) in sofrel; fold (so_func_related mfin e so) in sofrel.
        unfold S.ADC_step; unfold _get_st; unfold bind_s;
        unfold bind; simpl.
        rewrite cp_b; rewrite sd; simpl.
        apply (hasSPSR_false e m7 Events.E0 m7 v3
          (Arm6_State.set_reg s d
            (add (add (Arm6_State.reg_content s n) so)
              (Arm6_State.cpsr s) [Cbit]))
          ) in spsr_b;
          [idtac |inv spsr_b].
        unfold if_CurrentModeHasSPSR. unfold block. unfold fold_left.
        unfold _get_bo. unfold bind_s. unfold next. unfold bind.
        simpl; unfold _Arm_State.set_reg.
        rewrite spsr_b; simpl.
        exact psrel. exact hasspsr. 
      (* ((S == 1) && (d == 15)) evaluates to false *)
      apply (S_set_and_is_pc_false e m6 Events.E0 m6 v2 sbit d) in sd_b;
        [idtac|exact sfrel|exact dfrel|exact sd].
      inv main_p;
      rename H5 into is_s, H8 into s_b, H9 into main_p, H4 into evs;
          simpl in s_b; 
          apply no_effect_is_S_set in is_s;
          inversion is_s;
          rewrite H in * |- *;
          clear H is_s; rename H0 into is_s(* m6=m7*);
          apply Events.Eapp_E0_inv in evs; destruct evs; subst.      
        (* S == 1 evaluates to true *)
        inv main_p ;[idtac | nod];
        rename H4 into nf, H7 into main_p, H3 into evs;
        apply Events.Eapp_E0_inv in evs; destruct evs; subst.

        apply (S_is_set e m7 Events.E0 m7 v3 sbit) in s_b;
          [idtac|exact sfrel|exact is_s].

        inv nf; rename H2 into nf;
        pose (s0 :=  Arm6_State.set_reg s d
                       (add (add (Arm6_State.reg_content s n) so)
                          (Arm6_State.cpsr s) [Cbit]));
        fold s0 in psrel;
        eapply (same_nflag_assgnt e m7 nil (Util.zne d 15)
          s0 d Events.E0 m8 v4)
          in psrel;
          [idtac | exact dfrel | exact nf].

        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (nf_params_not_changed m7 e v4 m8 S) in sfrel;
          [idtac | exact nf];
        fold (bit_proj m8 e S) in sfrel; fold (sbit_func_related m8 e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert_fixed.cond) in cfrel;
          [idtac | exact nf];
        fold (cond_proj m8 e) in cfrel; fold (cond_func_related m8 e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert_fixed.d) in dfrel;
          [idtac | exact nf];
        fold (reg_proj m8 e adc_compcert_fixed.d) in dfrel; fold (d_func_related m8 e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert_fixed.n) in nfrel;
          [idtac | exact nf]; 
        fold (reg_proj m8 e adc_compcert_fixed.n) in nfrel; fold (n_func_related m8 e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (nf_params_not_changed m7 e v4 m8 shifter_operand) in sofrel;
          [clear nf | exact nf];
        fold (bits_proj m8 e shifter_operand) in sofrel; fold (so_func_related m8 e so) in sofrel.
        inv main_p ;[idtac | nod];
        rename H4 into zf, H7 into main_p, H3 into evs;
        apply Events.Eapp_E0_inv in evs; destruct evs; subst.

        inv zf; rename H2 into zf;
        pose (s1 := Arm6_State.set_cpsr_bit s0 Nbit
                       (Arm6_State.reg_content s0 d) [n31]);
        revert psrel; fold s1; intro psrel;
        eapply (same_zflag_assgnt e m8 nil (Util.zne d 15)
          s1
          d Events.E0 m9 v5) in psrel;
        [idtac| exact dfrel | exact zf].
        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (zf_params_not_changed m8 e v5 m9 S) in sfrel;
          [idtac | exact zf];
        fold (bit_proj m9 e S) in sfrel; fold (sbit_func_related m9 e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert_fixed.cond) in cfrel;
          [idtac | exact zf];
        fold (cond_proj m9 e) in cfrel; fold (cond_func_related m9 e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert_fixed.d) in dfrel;
          [idtac | exact zf];
        fold (reg_proj m9 e adc_compcert_fixed.d) in dfrel; fold (d_func_related m9 e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert_fixed.n) in nfrel;
          [idtac | exact zf]; 
        fold (reg_proj m9 e adc_compcert_fixed.n) in nfrel; fold (n_func_related m9 e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (zf_params_not_changed m8 e v5 m9 shifter_operand) in sofrel;
          [clear zf | exact zf];
        fold (bits_proj m9 e shifter_operand) in sofrel; fold (so_func_related m9 e so) in sofrel.
        inv main_p ;[idtac | nod];
        rename H4 into cf, H7 into vf, H3 into evs;
        apply Events.Eapp_E0_inv in evs; destruct evs; subst.
        inv cf; rename H2 into cf;
        pose (s2 := Arm6_State.set_cpsr_bit s1 Zbit
                       (if Util.zeq (Arm6_State.reg_content s1 d) 0
                        then repr 1
                        else repr 0));
        revert psrel; fold s2; intro psrel;
        eapply (same_cflag_assgnt m9 e nil (Util.zne d 15)
          s s2
          n so Events.E0 m10 v6) in psrel;
        [idtac| exact nfrel | exact sofrel| exact cf]. 
        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (cf_params_not_changed m9 e v6 m10 S) in sfrel;
          [idtac | exact cf];
        fold (bit_proj m10 e S) in sfrel; fold (sbit_func_related m10 e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert_fixed.cond) in cfrel;
          [idtac | exact cf];
        fold (cond_proj m10 e) in cfrel; fold (cond_func_related m10 e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert_fixed.d) in dfrel;
          [idtac | exact cf];
        fold (reg_proj m10 e adc_compcert_fixed.d) in dfrel; fold (d_func_related m10 e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert_fixed.n) in nfrel;
          [idtac | exact cf]; 
        fold (reg_proj m10 e adc_compcert_fixed.n) in nfrel; fold (n_func_related m10 e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (cf_params_not_changed m9 e v6 m10 shifter_operand) in sofrel;
          [clear cf | exact cf];
        fold (bits_proj m10 e shifter_operand) in sofrel; fold (so_func_related m10 e so) in sofrel.

        unfold st in psrel.
        inv vf; rename H2 into vf;
        pose (s3 := Arm6_State.set_cpsr_bit s2 Cbit
                       (Arm6_Functions.CarryFrom_add3
                         (Arm6_State.reg_content s n) so
                         (Arm6_State.cpsr s2) [Cbit]));
        revert psrel; fold s3; intro psrel;
        eapply (same_vflag_assgnt m10 e nil (Util.zne d 15)
          s s3
          n so Events.E0 mfin v7) in psrel;
        [clear vf| exact nfrel | exact sofrel| exact vf].

        unfold S.ADC_step. unfold _get_st. unfold bind_s; unfold bind; simpl.
        rewrite cp_b. simpl. 
        unfold block. unfold fold_left at 1. unfold next. 
        unfold bind at 1 2. unfold _get_bo at 1. 
        unfold bind_s at 1. unfold bind at 1. unfold bind at 1. 
        unfold set_reg. simpl; unfold _Arm_State.set_reg. 
        fold s0. 
        rewrite sd_b; rewrite s_b; simpl.
        (* Nflag *)
        unfold bind at 5. unfold _get_bo at 2. unfold bind_s at 1. 
        unfold bind at 5. unfold bind at 5.
        simpl; unfold _Arm_State.set_cpsr_bit at 1. 
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        unfold _set_bo at 1.  simpl. unfold ok_semstate.
        
        (* Zflag *)
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
        (* Cflag *)
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
        (* Vflag *)
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
        unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
        simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
        unfold bind at 4. unfold loc at 1. unfold bo at 1. unfold bo at 3.
        unfold st at 1. unfold st at 3.
        unfold bind at 3. unfold loc at 1. unfold bo at 1. unfold bo at 5.
        unfold st at 1. unfold st at 5.
        unfold bind at 2. unfold loc at 1. unfold bo at 1. unfold bo at 9.
        unfold st at 1. unfold st at 9.
        
        unfold bind at 1. unfold _get_bo at 2. unfold bind_s at 1.
        unfold bind at 1. unfold bo at 1.
        unfold _set_bo at 1. unfold loc at 1. unfold st at 1.
        unfold ok_semstate.
        unfold _get_bo at 1. unfold bind_s at 1. unfold bind at 1.
        unfold loc at 1. unfold bo. unfold st at 1. unfold st.
        fold s1. fold s2. fold s3. unfold st in psrel.
        rewrite same_bool; rewrite same_bool; rewrite same_bool;
        rewrite same_bool; rewrite same_bool.
        exact psrel.

        (* S == 1 evaluates to false *)
        inv main_p.
        apply (S_not_set e mfin Events.E0 mfin v3 sbit) in s_b;
          [idtac|exact sfrel|exact is_s].
        unfold S.ADC_step; unfold _get_st; unfold bind_s; unfold bind; simpl.
        rewrite cp_b; rewrite sd_b; rewrite s_b; simpl.
        unfold block. unfold fold_left. unfold next.
        unfold bind at 3. simpl; unfold _Arm_State.set_reg.
        unfold _get_bo at 2. unfold bind_s at 1. unfold _set_bo at 1.
        unfold ok_semstate.
        unfold bind at 3. unfold loc at 1. unfold bo at 1.
        unfold st at 1.
        unfold _get_bo at 1. unfold bind_s at 1. unfold bind at 3.
        unfold bind at 2.
        unfold bind at 2. unfold _get_bo at 1. unfold bind_s at 1.
        unfold bind at 2. unfold _get_bo at 1. unfold bind_s at 1.
        unfold _set_bo at 1. unfold ok_semstate.
        unfold bind at 2.
        unfold bind at 1. unfold loc. unfold bo. unfold st. simpl.
        simpl. rewrite same_bool. exact psrel. (*exact condpass0. exact condpass0.*)

    (* ConditionPassed(&proc->cpsr, cond) evaluates to false *)
    inv main_p.
    unfold S.ADC_step; unfold _get_st; unfold bind_s; unfold bind; simpl.
    rewrite (condpass_false m0 m1 e mfin Events.E0 mfin v1);
      [simpl;exact psrel |exact al| exact condpass0 |exact cp_b].
Qed.

