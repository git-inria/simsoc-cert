Require Import Globalenvs Memory.
Require Import Csyntax Csem Cstrategy Coqlib Integers Values Maps Errors. 
Require Import Arm6_State Arm6_Proc Arm6_SCC Bitvec Arm6.
Require Import adc_compcert.
Require Import projection. 

Require Import Arm6_Simul.
Import I.
Import Arm6_Functions.Semantics.

(* Functional relation between the C memory module which contains the other ADC parameters, 
   and the COQ specification of ADC parameters *)
Definition sbit_func_related (m:Mem.mem) (e:env) (sbit:bool):Prop:=
  bit_proj m e S = sbit.

Definition cond_func_related (m:Mem.mem) (e:env) (cond:opcode):Prop:=
  cond_proj m e = cond.

Definition d_func_related (m:Mem.mem) (e:env) (d:regnum):Prop:=
  reg_proj m e adc_compcert.d = d.

Definition n_func_related (m:Mem.mem) (e:env) (n:regnum):Prop:=
  reg_proj m e adc_compcert.n = n.

Definition so_func_related (m:Mem.mem) (e:env) (so:word):Prop:=
  bits_proj m e shifter_operand = so.

(* Human readable renaming of [p], which is generated by the Coq printer *)
Definition prog_adc := adc_compcert.p.

(* The assignment of old_Rn has a normal outcome *)
Lemma normal_outcome_for_assgnt: 
  forall a1 a2 ge t ev m e m' out,
  exec_stmt ge e m (Sdo (Eassign a1 a2 t)) ev m' out ->
  out = Out_normal.
Proof.
intros until out. intros exst. 
inv exst. reflexivity.
Qed.

Implicit Arguments normal_outcome_for_assgnt [a1 a2 ge t ev m e m' out].

Ltac noa :=
  match goal with
    [He: exec_stmt _ _ _ (Sdo (Eassign _ _ _)) _ _ ?out,
     Hd: ?out <> Out_normal |- _ ] =>
       case Hd; 
       apply (normal_outcome_for_assgnt He) end.

(* Any Sdo has a normal outcome*)
Lemma normal_outcome_for_do:
  forall exp ge t m e m' out,
    exec_stmt ge e m (Sdo exp) t m' out ->
    out = Out_normal.
Proof.
  intros until out. intros exst.
  inv exst. reflexivity.
Qed.

Implicit Arguments normal_outcome_for_do [exp ge t m e m' out].

Ltac nod :=
  match goal with
    [He: exec_stmt _ _ _ (Sdo _) _ _ ?out,
     Hd: ?out <> Out_normal |- _ ] =>
       case Hd; 
       apply (normal_outcome_for_do He) end.  



(* Return the memory model which only relates to this ident *)
Parameter of_mem : AST.ident -> Mem.mem -> Mem.mem.

(*exp get_bit*)
Print fun_internal_ADC.

Definition reg_id id :=
  Ecall (Evalof (Evar reg T2) T2)
  (Econs (Evalof (Evar proc T3) T3)
    (Econs 
      (Evalof (Evar id T4) T4) Enil)) T1.

Definition get_rd_bit31 :=
  Ecall (Evalof (Evar get_bit T17) T17)
  (Econs (reg_id d)
    (Econs (Eval (Vint (repr 31)) T9)
      Enil)) T10.

Lemma same_reg_d :
  forall e m t m' a' l b st d,
    proc_state_related m e (Ok tt (mk_semstate l b st)) ->
    d_func_related m e d ->    
    eval_expr (Genv.globalenv prog_adc) e m RV 
              (reg_id adc_compcert.d) t m' a' ->
    a'= (Eval (Vint (Arm6_State.reg_content st d)) T1).
Admitted.

Set Implicit Arguments.

Lemma alloc_diff_block :
  forall m e e' m' x y b_x tx b_y ty,
    alloc_variables e m ((x,tx)::(y,ty)::nil) e' m'->
    list_norepet (x::y::nil) ->
    e' ! x = Some (b_x, tx) ->
    e' ! y = Some (b_y, ty) ->
    b_x <> b_y.
Proof.
  intros until ty. intros av norepet getx gety.
  inv av. inv H7. inv H9.
  apply Mem.valid_new_block in H6.
  unfold Mem.valid_block in H6.
  apply Mem.alloc_result in H8.
  rewrite <- H8 in H6; clear H8.
(* SearchPattern (_ < _ -> _ <> _). *)
  apply Zlt_not_eq in H6.
  assert (findy: (PTree.set y (b0, ty) (PTree.set x (b1, tx) e)) ! y =
                  Some (b0, ty)).
  apply PTree.gss. rewrite findy in gety. inversion gety.

  assert (findx: (PTree.set y (b0, ty) (PTree.set x (b1, tx) e)) ! x =
                  (PTree.set x (b1, tx) e) ! x).
  apply PTree.gso.
  inv norepet. unfold In in H2. intro exy. apply H2. left. symmetry. exact exy.

(*info intuition.*)

  rewrite findx in getx.
  rewrite PTree.gss in getx. inversion getx.
  rewrite <- H0. rewrite <- H1.
  exact H6.
Qed.

Lemma lt_block :
  forall m1 ofs1 b1 m2 ofs2 b2 m3,
    Mem.alloc m1 0 ofs1 = (m2, b1) ->
    Mem.alloc m2 0 ofs2 = (m3, b2) ->
    b1 < b2.
Proof.
  intros until m3. intros alc1 alc2.
  apply Mem.valid_new_block in alc1. unfold Mem.valid_block in alc1.
  apply Mem.alloc_result in alc2. rewrite <- alc2 in alc1.
  exact alc1.
Qed.


Ltac blocks_lt b1 b2 :=
  match goal with [alc1: Mem.alloc ?m1 ?l1 ?h1 = (?m2, b1) |- ?c1 ]=>
    match goal with
      |[alc2: Mem.alloc m2 ?l2 ?h2 = (?m3, b2) |- ?c ] =>
        apply lt_block with m1 h1 b1 m2 h2 b2 m3 in alc1;
          [idtac|exact alc2]
      |[alc2: Mem.alloc ?mx ?lx ?hx = (?my, ?bx) |- ?c ] =>
        apply lt_block with m1 h1 b1 mx hx bx my in alc1;
          [blocks_lt bx b2|exact alc2]
    end
  end.

Ltac blocks_lt' b1 b2 :=
  match goal with
    |[lt1: b1 < b2 |- ?c] => idtac
    |[lt1: b1 < ?bx |- ?c] =>
      match goal with
        |[lt2: bx < b2 |- ?c] => 
          apply (Zlt_trans b1) in lt2;
            [clear lt1|exact lt1]
        |[lt2: bx <?bxx |-?c]=>
          try apply (Zlt_trans b1) in lt2;
            [clear lt1;blocks_lt' b1 b2|exact lt1]
      end
  end.

Ltac blocks_neq b1 b2 :=
  match goal with
    |[lt1: b1 < b2 |- ?c] => apply Zlt_not_eq in lt1
    |[lt1: b1 < ?bx |- ?c] =>
      match goal with
        |[lt2: bx < b2 |- ?c] => 
          apply (Zlt_trans b1) in lt2;
            [clear lt1;apply Zlt_not_eq in lt2|exact lt1]
        |[lt2: bx <?bxx |-?c]=>
          try apply (Zlt_trans b1) in lt2;
            [clear lt1;blocks_neq b1 b2|exact lt1]
      end
  end.

Ltac diff_blk b1 b2:=
  blocks_lt b1 b2; blocks_neq b1 b2.

Lemma diff_block :
  forall m1 ofs1 b1 m2 ofs2 b2 m3,
    Mem.alloc m1 0 ofs1 = (m2, b1) ->
    Mem.alloc m2 0 ofs2 = (m3, b2) ->
    b1 <> b2.
Proof.
  intros until m3. intros alc1 alc2.
  apply Mem.valid_new_block in alc1. unfold Mem.valid_block in alc1.
  apply Mem.alloc_result in alc2. rewrite <- alc2 in alc1.
  apply Zlt_not_eq in alc1.
  exact alc1.
Qed.

Set Printing Depth 30.
(*
Lemma and_zdiv_1:
  forall (x:word) (n:Z),
    0 < n < Z_of_nat wordsize ->
    (repr n) = x -> and (repr n) x / n = 1.
Proof.
  intros. rewrite <- H0. SearchAbout and. rewrite and_idem.
  SearchAbout Zdiv. 
*)
Lemma same_getbit :
  forall x n ,
    0 < n < Z_of_nat wordsize ->
    sign_ext 8 (and (shru x (repr n)) (repr 1)) = x [nat_of_Z n].
Proof.
(*  intros.
  assert (0 < 8 < Z_of_nat wordsize).
  simpl. omega.
  apply zero_ext_and with (x := (and (shru x (repr n)) (repr 1))) in H0.
  rewrite H0.  
  unfold bit. unfold bits. unfold bits_val.
  unfold masks. (*SearchAbout minus. *)
  rewrite minus_diag. (*Print masks_aux.*)
  simpl masks_aux. 
  (*SearchAbout repr.*)
  rewrite shru_div_two_p.
*)
(*
  induction n. 
  simpl nat_of_Z. 
  unfold masks. simpl masks_aux.
  rewrite two_power_nat_O.
  SearchAbout (Zdiv).
  rewrite Zdiv_1_r.
  (*lemma on 'repr' apply eqm_samerepr. apply eqm_refl2.*)
  SearchAbout two_p.
  assert (8 = Z_of_nat 8).
  simpl; reflexivity. rewrite H0.
  rewrite <- two_power_nat_two_p.
  rewrite Word.shru_zero.
  SearchAbout and.
  admit.
  admit.
  unfold nat_of_Z.
  unfold masks. simpl masks_aux.
  rewrite two_power_nat_O.
  rewrite Zdiv_1_r.
  assert (8 = Z_of_nat 8).
  simpl; reflexivity. rewrite H0.
  rewrite <- two_power_nat_two_p.
  SearchAbout Zneg.
*)
Admitted.

(* expirement on how to avoid using inversion *)
(*
Ltac gen_inv_S y :=
 pattern y; 
 match goal with [ |- ?concl _ ] => 
   change (match S y with S y => concl y | _ => True end) end;
 cbv beta.
*)

(* simplify the inversion on alloc_variables and bind_parameters definition *)
Ltac inv_alloc_vars e' :=
  let ex :=fresh "e" in
  let mx :=fresh "m" in
  let idx :=fresh "id" in
  let tyx :=fresh "ty" in
  let varsx :=fresh "vars" in
  let m1x :=fresh "m1" in
  let b1x :=fresh "b1" in
  let m2x :=fresh "m2" in
  let e2x :=fresh "e2" in
  let alc :=fresh "alc" in
  let av' := fresh "av'" in
  match goal with 
    [av: alloc_variables ?e ?m0 ?lst e' ?m0' |- ?c] => 
    inversion av as [ex mx|ex mx idx tyx varsx m1x b1x m2x e2x alc av'];
    subst;try clear av;
    (inv_alloc_vars e'||idtac)
  end.

Ltac inv_bind_params m' :=
  let ex :=fresh "e" in
  let mx :=fresh "m" in
  let idx :=fresh "id" in
  let tyx :=fresh "ty" in
  let paramsx :=fresh "params" in
  let v1x :=fresh "v1" in
  let vlx :=fresh "vl" in
  let bx :=fresh "b" in
  let m1x :=fresh "m1" in
  let m2x :=fresh "m2" in
  let eget :=fresh "eget" in
  let str :=fresh "str" in
  let bp' := fresh "bp'" in
  let Heq := fresh "Heq" in
  match goal with
    [bp: bind_parameters ?e ?m ?lst ?vlst m' |- ?c] =>
    inversion bp as 
      [ex mx Heq
        |ex mx idx tyx paramsx v1x vlx bx m1x m2x eget str bp'];
    try clear bp;subst;try simpl in eget;
    (inv_bind_params m'|| idtac)
  end.

Ltac rrw_block :=
  let Heq := fresh "Heq" in
  match goal with [eq:Some ?l = Some (?b,?t)|-?c] => 
    injection eq;intro Heq;rewrite<-Heq in *;clear Heq eq b end.

(* The loaded value from block b is not changed between m1, m2.
   From m1 to m2, we consider all the storage in memory. 
   If there is no store on block b, then the value in b is not changed *)
Ltac val_not_changed_str ck b o m m' :=
  match goal with
    |[str1: Mem.store ?ck1 m b ?ofs1 ?v1 = Some ?m2 |-?c]=>idtac
    |[str1: Mem.store ?ck1 m ?b1 ?ofs1 ?v1 = Some m' |-?c]=>
      generalize str1;
      apply Mem.load_store_other with ck1 m b1 ofs1 v1 m' ck b o in str1;
        [idtac|left;diff_blk b b1;assumption]
    |[str1: Mem.store ?ck1 m ?b1 ?ofs1 ?v1 = Some ?m2 |-?c]=>
      match goal with
        |[str2: Mem.store ?ck2 m2 ?b2 ?ofs2 ?v2 = Some ?m3|-?c]=>
          generalize str1;
          apply Mem.load_store_other with ck1 m b1 ofs1 v1 m2 ck b o in str1;
            [idtac|left;diff_blk b b1;assumption];
          val_not_changed_str ck b o m2 m'
      end
  end.

Ltac case_I h := case h; try (intros; exact I); clear h.

Ltac case_h h := case h; clear h; try contradiction.

Ltac rew_clean eq :=
  match type of eq with ?l = ?r => rewrite eq in *; clear eq l end.

Ltac and_eq_subst ae :=
  repeat (rew_clean ae) ||
         (let feq := fresh "eq" in destruct ae as [feq ae];
          rew_clean feq).

Ltac inv_end ev mm mm' :=
   unfold ev, mm, mm' in *; clear ev mm mm'; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_ecall_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env arg_m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?c] =>
    pose (e := Ecall a1 a2 a3); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert 
      (em : match e with 
                      |Ecall a b c =>
                        (a=a1)/\(b=a2)/\(c=a3)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                      |_=> False
                    end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.

Ltac inv_ecall arg_m t1 m2 rf' t2 m3 rargs' 
         vf vargs0 targs tres fd t3 vres H H0 H1 H2 H3 H4 H5 H6 :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_ecall_begin arg_m ev mm mm'; 
  intros e0 m1 rf rargs ty t1 m2 rf' t2 m3 rargs' 
         vf vargs0 targs tres fd t3 m4 vres H H0 H1 H2 H3 H4 H5 H6;
  inv_end ev mm mm'.

Ltac inv_evalof_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env arg_m _ (Evalof ?a1 ?a2) _ ?m' _ |- ?c ] =>
    pose (e := Evalof a1 a2); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert 
      (em : match e with 
                    |Evalof a b => 
                      (a=a1)/\(b=a2)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                    |_ => False
                  end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.

Ltac inv_evalof arg_m t0 m'0 a' H :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_evalof_begin arg_m ev mm mm'; 
  intros e0 m1 a t0 m'0 a' ty H;
  inv_end ev mm mm'.

Ltac inv_evar_begin arg_m ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h: eval_expr _ ?env arg_m _ (Evar ?a1 ?a2) _ ?m' _ |- ?c] =>
    pose (e := Evar a1 a2); 
    pose (ev:=env); pose (mm:=arg_m); pose (mm':=m');
    assert
      (em: match e with
                   |Evar a b => 
                     (a=a1)/\(b=a2)/\(env=ev)/\(arg_m=mm)/\(m'=mm')
                   |_ => False
                 end)
      by repeat (split||reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.
  
Ltac inv_evar arg_m :=
  let ev:=fresh "ev" in 
  let mm:=fresh "mm" in 
  let mm':=fresh "mm'" in
  inv_evar_begin arg_m ev mm mm';
  intros e0 m1 x ty;
  inv_end ev mm mm'. 

Ltac inv_evalof_simplrv_begin v :=
  match goal with [h: eval_simple_rvalue _ _ _ (Evalof ?a1 ?a2) v |- ?c] =>
    let e := fresh "expr" in
    pose (e := Evalof a1 a2);
    assert
      (rm: match e with
                   |Evalof a b =>(a = a1) /\ (b = a2)
                   |_=>False
                 end)
      by repeat  (split||reflexivity);
    fold e in h;
    revert rm;
    case_h h;
    clear e
  end.

Ltac inv_evalof_simplrv_end :=
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_evalof_simplrv v b0 ofs v0 H H0 H1 :=
  inv_evalof_simplrv_begin v;
  intros b0 ofs l0 ty v0 H H0 H1;
  inv_evalof_simplrv_end. 

Ltac inv_av_cons_begin arg_m ev :=
  let lst := fresh "lst" in
  match goal with [av: alloc_variables ?env arg_m ((?id,?ty) ::?t) ?a3 ?a4 |- ?c] => 
    pose (lst := ((id,ty)::t)); pose (ev:=env);
    change (alloc_variables ev arg_m lst a3 a4) in av;
    assert
      (lm: match lst with
                    |(a,b)::c=>(a=id)/\(b=ty)/\(c=t)/\(ev=env)
                    |_=>False
                  end)
      by repeat (split||reflexivity);
    revert lm;
    case_h av;
    clear lst
  end.

Ltac inv_av_cons_end ev :=
   unfold ev in *; clear ev; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).  

Ltac inv_av_cons arg_m m m1 b1 m4 e2 H H0:=
  let ev:=fresh "ev" in 
  inv_av_cons_begin arg_m ev;
  intros e0 m id0 ty vars m1 b1 m4 e2 H H0;
  inv_av_cons_end ev.

Ltac inv_av_nil_begin arg_m lnil ev ev' :=  
  match goal with [av: alloc_variables ?env arg_m ?lst ?env' ?a4 |- ?c] =>
    pose (lnil:=lst); pose (ev:=env); pose (ev':=env');
    change (alloc_variables ev arg_m lnil ev' a4) in av;
    assert (lm:match lnil with 
                        |nil =>(nil = lst)/\(ev=env)/\(ev'=env')
                        |_ =>False end) 
      by repeat (split||reflexivity);
    revert lm;
    case_h av    
  end.

Ltac inv_av_nil_end lnil ev ev' :=
   unfold lnil, ev, ev' in *; clear lnil ev ev'; 
   let ae := fresh "ae" in (intro ae; and_eq_subst ae).

Ltac inv_av_nil arg_m e0 m :=
  let lnil:=fresh "lnil" in 
  let ev:=fresh "ev" in 
  let ev':=fresh "ev'" in 
  inv_av_nil_begin arg_m lnil ev ev';
  intros e0 m;
  inv_av_nil_end lnil ev ev'.  

(*
Definition inv_expr_ecall e m ex m' (ex':expr):=
  match ex with
    |Ecall a b c => 
      forall (X:Prop), 
      (forall g t1 m1 rf' t2 m2 rargs' vf vargs targs tres fd t3 vres,
      eval_expr g e m RV a t1 m1 rf' -> 
      eval_exprlist g e m1 b t2 m2 rargs' ->
      eval_simple_rvalue g e m2 rf' vf ->
      eval_simple_list g e m2 rargs' targs vargs ->
      typeof a = Tfunction targs tres ->
      Genv.find_funct g vf = Some fd ->
      type_of_fundef fd = Tfunction targs tres ->
      eval_funcall g m2 fd vargs t3 m' vres -> X) -> X
    |_=> True
  end.
*)

(* Auxiliary functions for inversion on type eval_expr *)
(* Constructor eval_call *)

Definition inv_expr_ecall' g e m ex m' ex':=
  match ex with
    |Ecall a b c as ecall =>
      forall (X:expr -> Prop),
      (forall rf t1 m1 rf' t2 m2 rargs' vf vargs targs tres fd t3 vres,
      eval_expr g e m RV a t1 m1 rf' -> 
      eval_exprlist g e m1 b t2 m2 rargs' ->
      eval_simple_rvalue g e m2 rf' vf ->
      eval_simple_list g e m2 rargs' targs vargs ->
      classify_fun (typeof rf) = fun_case_f targs tres->
      (*typeof a = Tfunction targs tres ->*)
      Genv.find_funct g vf = Some fd ->
      type_of_fundef fd = Tfunction targs tres ->
      eval_funcall g m2 fd vargs t3 m' vres -> 
      X (Eval vres (typeof ecall))) -> X ex'
    |_=> True
  end.

(* Constructor eval_valof *)
Definition inv_expr_valof g e m ex m' ex' :=
  match ex with
    |Evalof b c as evalof=>
      forall (X:expr->Prop),
        (forall t a',
          eval_expr g e m LV b t m' a'->X (Evalof a' (typeof evalof)))->
          X ex'
    |_=>True
  end.

(* General inversion tactic on eval_expr from m to m' *)
Ltac inv_eval_expr m m' :=
  let f:=fresh "f" in
  let nexp:=fresh "nexp" in
  let a_:=fresh "a" in
  let a'_:=fresh "a'" in
  (*ev_funcall*)
  let rf_:=fresh "rf" in
  let t1_:=fresh "t" in
  let t2_:=fresh "t" in
  let t3_:=fresh "t" in
  let m1_:=fresh "m" in
  let m2_:=fresh "m" in
  let rf'_:= fresh "rf'" in
  let rargs'_:=fresh "rargs'" in
  let vf_:=fresh "vf" in
  let vargs_:=fresh "vargs" in
  let targs_:=fresh "targs" in
  let tres_:=fresh "tres" in
  let fd_:=fresh "fd" in
  let vres_:=fresh "vres" in
  let ty_:=fresh "ty" in
  let ev_ex:=fresh "ev_ex" in
  let ev_elst:=fresh "ev_eslst" in
  let esr1:=fresh "esr" in
  let esr2:=fresh "esr" in
  let Heqcf:=fresh "Heqcf" in
  let eslst:=fresh "eslst" in
  let Heqff:=fresh "Heqff" in
  let Heqtf:=fresh "Heqtf" in
  let ev_funcall:=fresh "ev_funcall" in
  match goal with
    |[ee:eval_expr ?ge ?e m RV (Econdition ?a1 ?a2 ?a3 ?ty) ?t ?m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1: eval_expr ge e m RV a1 ?t1 ?mcond ?a1'|-?cl1]=>
          inv_eval_expr m mcond
      end
    |[ee:eval_expr ?ge ?e m RV (Eval ?v ?ty) ?et m' ?a'|-?cl]=>
      inv ee
    |[ee:eval_expr ?ge ?e m LV (Evar ?x ?ty) ?et m' ?a'|-?cl]=>
      inv ee
    |[ee:eval_expr ?ge ?e m RV (Ebinop ?op ?a1 ?a2 ?ty) ?t m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1:eval_expr ?ge ?e m ?k a1 ?t1 ?mbo ?a1'|-?cl1]=>
          inv_eval_expr m mbo;inv_eval_expr mbo m'
      end
    |[ee:eval_expr ?ge ?e m RV (Evalof ?a ?ty) ?t m' ?a'|-?cl]=>
      generalize
        (match ee in (eval_expr _ e m _ ex _ m' ex')
           return inv_expr_valof (Genv.globalenv prog_adc) e m ex m' ex' with
           |eval_valof _ _ a t _ a' ty H1 =>
             (fun X k => k t a' H1)
           |_=> I
         end);clear ee;
        intro k; red in k;simpl in k;
        pose(nexp:=a');change a' with nexp in k; 
          match goal with
            |[es:context c [a']|-?cl]=>revert es
            |_=>idtac
          end;
          unfold nexp in k;clear nexp;apply k;clear k;
          intros t1_ a_;intro ev_ex;intro esr1;
      (*inv ee;*)inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m LV (Efield ?a ?f ?ty) ?t m' ?a'|-?cl]=>
      inv ee;inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m LV (Ederef ?a ?ty) ?t m' ?a'|-?cl]=>
      inv ee;inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m RV (Eaddrof ?a ?ty) ?t m' ?a'|-?cl]=>
      inv ee;inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m RV (Eunop ?op ?a ?ty) ?t m' ?a'|-?cl]=>
      inv ee;inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m RV (Ecast ?a ?ty) ?t m' ?a'|-?cl]=>
      inv ee;inv_eval_expr m m'
    |[ee:eval_expr ?ge ?e m RV (Esizeof ?ty' ?ty) ?t m ?a'|-?cl]=>
      inv ee
    |[ee:eval_expr ?ge ?e m RV (Eassign ?l ?r ?ty) ?t m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1:eval_expr ge e m LV l ?t1 ?masgn1 ?l'|-?cl]=>
          inv_eval_expr m masgn1;
          match goal with
            |[ee2:eval_expr ge e masgn1 RV r ?t2 ?masgn2 ?r'|-?cl]=>
              inv_eval_expr masgn1 masgn2
          end
      end
    |[ee:eval_expr ?ge ?e m RV (Eassignop ?op ?l ?r ?tyres ?ty) ?t m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1:eval_expr ge e m LV l ?t1 ?masgnop1 ?l'|-?cl]=>
          inv_eval_expr m masgnop1;
          match goal with
            |[ee2:eval_expr ge e masgnop1 RV r ?t2 ?masgnop2 ?r'|-?cl]=>
              inv_eval_expr masgnop1 masgnop2
          end
      end
    |[ee:eval_expr ?ge ?e m RV (Epostincr ?id ?l ?ty) ?t m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1:eval_expr ge e m LV l t ?mpi ?l'|-?cl]=>
          inv_eval_expr m mpi
      end
    |[ee:eval_expr ?ge ?e m RV (Ecomma ?r1 ?r2 ?ty) ?t m' ?a'|-?cl]=>
      inv ee;
      match goal with
        |[ee1:eval_expr ge e m RV r1 ?t1 ?mcom ?r1'|-?cl]=>
          inv_eval_expr m mcom; inv_eval_expr mcom m'
      end
    |[ee:eval_expr ?ge ?e m RV (Ecall ?rf ?rargs ?ty) ?t m' ?a'|-?cl]=>
      generalize 
        (match ee in (eval_expr _ e m _ ex _ m' ex')
           return inv_expr_ecall' (Genv.globalenv prog_adc) e m ex m' ex' with
           |eval_call _ _ rf rargs typ t1 m1 rf' t2 m2 rargs' vf vargs
             targs tres fd t3 _ vres H1 H2 H3 H4 H5 H6 H7 H8 =>
             (fun X k => k rf t1 m1 rf' t2 m2 rargs' vf vargs 
               targs tres fd t3 vres H1 H2 H3 H4 H5 H6 H7 H8 )
           |_=> I
         end);clear ee;
        intro k;red in k;simpl in k;
        pose(nexp:=a');fold nexp in k;
        match goal with
          |[es:context [a']|-?cl]=>revert es
        end;
        unfold nexp in k;clear nexp;apply k;clear k;
        intros rf_ t1_ m1_ rf'_ t2_ m2_ rargs'_ vf_ vargs_ targs_ tres_ fd_ t3_ 
          vres_;
        intros ev_ex ev_elst esr1 eslst Heqcf Heqff Heqtf 
          ev_funcall esr2;
      match goal with
        |[ee1:eval_expr ge e m RV rf ?t1 ?mc1 ?rf'|-?cl]=>
          inv_eval_expr m mc1;
          match goal with
            |[eel:eval_exprlist ge e mc1 ?rargs ?t2 ?mc2 ?rargs'|-?cl]=>
              inv_eval_expr mc1 mc2
          end
      end
    |[eel:eval_exprlist ?ge ?e m (Econs ?a1 ?al) ?t m' ?rargs'|-?cl]=>
      inv eel;
      match goal with
        |[eel1:eval_expr ge e m RV a1 ?t1 ?ml1 ?a1'|-?cl]=>
          inv_eval_expr m ml1; inv_eval_expr ml1 m'
      end
    |[eel:eval_exprlist ?ge ?e m Enil ?t m' ?al'|-?cl]=>
      inv eel
    |_=> pose(f:=0)
  end.


Lemma same_get_reg' :
  forall e m0 m0' vargs m l b s d t m' v,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    proc_state_related m e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m get_rd_bit31  t m' v->
    v = Vint ((Arm6_State.reg_content s d) [n31]).
Proof.
  intros until v. intros av bp psrel dfrel get_bit.
  
  inversion get_bit as [env m1 gb t1 m1' gb' v1 gb_expr ev_rv Heqenv Heqm
    Heqexp Heqt Heqm' Heqv]; clear get_bit; subst.

  unfold get_rd_bit31 in gb_expr.


(*  revert ev_rv.
*)

(** new thought *)
(** Using impredicative encoding in inversion tactic *)
generalize 
  (match gb_expr in (eval_expr _ e m _ ex _ m' ex')
  return inv_expr_ecall' (Genv.globalenv prog_adc) e m ex m' ex' with
     |eval_call _ _ rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs
                      targs tres fd t3 _ vres H1 H2 H3 H4 H5 H6 H7 H8 =>
       (fun X k => k rf t1 m1 rf' t2 m2 rargs' vf vargs 
      targs tres fd t3 vres H1 H2 H3 H4 H5 H6 H7 H8 )
     |_=> I
   end). clear gb_expr.
intro k. red in k. simpl in k. revert ev_rv. apply k. clear k. 
intros until vres. 
intros gb_expr ev_explst ev_rv1 ev_simlst Heqty_gb Heqff Heqtyfd ev_funcall. 
intro ev_rv.

generalize 
  (match gb_expr in (eval_expr _ e m _ ex _ m' ex')
     return inv_expr_valof (Genv.globalenv prog_adc) e m ex m' ex' with
     |eval_valof _ _ a t _ a' ty H1 =>
       (fun X k => k t a' H1)
     |_=> I
   end). clear gb_expr.
intro k. red in k. simpl in k. revert ev_rv1. apply k. clear k.
intros until a'. intros gb_expr. intro ev_rv1.


(** Using impredicative encoding, 
   but without considering the output of expression evaluation *)
(*
generalize 
  (match gb_expr in (eval_expr _ e m _ ex _ m' ex')
  return inv_expr_ecall e m ex m' ex' with
     |eval_call e m rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs
                      targs tres fd t3 m3 vres H1 H2 H3 H4 H5 H6 H7 H8 =>
       (fun X k => k (Genv.globalenv prog_adc) t1 m1 rf' t2 m2 rargs' vf vargs 
                     targs tres fd t3 vres H1 H2 H3 H4 H5 H6 H7 H8)
     |_=> I
   end). clear gb_expr.
intro k. apply k. clear k.
*)

(** Without impredicative encoding *)
(* info 
  match goal with [h : eval_expr _ ?env ?m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?cl] =>
    let ex := fresh "expr_call" in
    pose (arg1 := a1);  
    pose (arg2 := a2);  
    pose (arg3 := a3);
    pose (ex := Ecall arg1 arg2 arg3);
    change (match ex with 
                      |Ecall a b c => cl
                      |_=> True
                    end);
    assert (ee : ex = Ecall arg1 arg2 arg3) by reflexivity; 
    revert ee;
    revert av bp psrel dfrel;
  
    change (Ecall a1 a2 a3) with ex in gb_expr;
    case gb_expr; try (intros; exact I); clear gb_expr e m t m' gb';
    intros e m rf rargs ty t1 m1 rf' t2 m2 rargs' vf vargs0 targs tres fd
      t3 m3 vres;
    intros gb_expr ev_exlst ev_simprv1 ev_simplst Heqtyrf Heqff Heqtyfd ev_funcall;
    intros av bp pstrl dfrel Heqexpr ev_simprv;
    injection Heqexpr; intros Heqty Heqrargs Heqrf;
    unfold arg1, arg2, arg3 in Heqty, Heqrargs, Heqrf; 
    clear arg1 arg2 arg3 Heqexpr expr_call;
    rewrite Heqty in ev_simprv;
    rewrite Heqrargs in ev_exlst;
    rewrite Heqrf in gb_expr, Heqtyrf;
    clear Heqty Heqrargs Heqrf
  end.
*)  

(* *********************************************************************)
(** old one *)
(** With extra equalities introduced in inversion tactic *)
(* 
Ltac inv_ecall_begin ev mm mm' :=
  let e := fresh "expr" in
  let em := fresh "expr_match" in
  match goal with [h : eval_expr _ ?env ?m _ (Ecall ?a1 ?a2 ?a3) _ ?m' _|- ?c] =>
    pose (e := Ecall a1 a2 a3); 
    pose (ev:=env); pose (mm:=m); pose (mm':=m');
    assert 
      (em : match e with 
                      |Ecall a b c =>
                        (a=a1)/\(b=a2)/\(c=a3)/\(env=ev)/\(m=mm)/\(m'=mm')
                      |_=> False
                    end)
      by repeat (split || reflexivity);
  fold e in h;
  revert em;
  case_h h;
  clear e
  end.
*)

(*
  inv_ecall m t1 m2 rf' t2 m3 rargs' vf vargs0 targs tres fd t3 vres
            gb_expr explst ev_rv1 ev_simlst H_ Heqfindfd Heqt16 ev_funcall. clear H_.
  intro ev_rv.
*)


(*
  (*harmless inversion: no ordering changes, no new hyp*)
  inversion ev_rv; subst; clear ev_rv.

  revert ev_rv1.
  inv_evalof m t0 m'0 a' H.
(*intro ev_rv1.

  revert ev_rv1.*)
  inv_evar m.
  intro ev_rv1.
  clear t0 a'.

  inv_evalof_simplrv vf b0 ofs v0 ev_simpl_lv Heqty Heqlvot.

  assert (globenv: e!get_bit=None).
    simpl in av.
    
    inv_av_cons m0 ma_proc m_proc b_proc m_proc' e_proc Heqma_proc av.
    inv_av_cons m_proc ma_s m_s b_s m_s' e_s Heqma_s av.
    inv_av_cons m_s ma_cond m_cond b_cond m_cond' e_cond Heqma_cond av.
    inv_av_cons m_cond ma_d m_d b_d m_d' e_d Heqma_d av.
    inv_av_cons m_d ma_n m_n b_n m_n' e_n Heqma_n av.
    inv_av_cons m_n ma_so m_so b_so m_so' e_so Heqma_so av.
    inv_av_cons m_so ma_on m_on b_on m_on' e_on Heqma_on av.

    inv_av_nil_begin m_on lnil ev ev'.
    intros.

    destruct lm as [feq ae]; clear feq.
    destruct ae as [feq ae]; rewrite feq in *; clear feq.
    rewrite <- ae in *; clear ae.

    
*)
    (*
    simpl; reflexivity.

  match goal with [_: eval_simple_lvalue _ _ _ (Evar ?a1 ?a2) _ _ |- ?c] =>
    assert
      (lv_match: match expr_evar with
                   |Evar a b =>(a = a1) /\ (b = a2)
                   |_=>False
                 end)
      by repeat  (split||reflexivity)
  end. 
  fold expr_evar in ev_lv.
  revert lv_match.

  case_h ev_lv.
    (*get_bit is in global environment *)
    intros until b1. intro locenv. intros.
    destruct lv_match as [eq1 eq2]; subst.
    rewrite locenv in globenv; discriminate.
    (*get_bit is in local environment *)
    intros until b1; intros _ Heqfindsymb _; intros.
    destruct lv_match as [eq1 eq2]; rewrite eq1 in *; clear eq1 eq2.*)

    (*match goal with [_:eval_exprlist _ _ _ (Econs ?a1 ?a2) _ _ _]*)
    
    
   
  

(* useful trick for later
  match goal with [_ : eval_expr _ _ _ _ ?interesting _ _ _ |- ?c ] => 
     let name := fresh e0 in 
     pose (name := interesting) end.
*)  

  (*revert gb_sim_rv.  
  generalize (refl_equal get_bit_reg).
  unfold get_bit_reg at 2.
  case gb_expr; clear gb_expr; try (intros; discriminate). 
  intros. injection H7. clear H7. intros; subst.*)


(*match goal with [ |- context c [Ecall ?a1 ?a2 ?a3]] => pattern a1, a2, a3 end.
    change 
      (match Ecall (Evalof (Evar get_bit T16) T16)
     (Econs (reg_id adc_compcert.d)
        (Econs (Eval (Vint (repr 31)) T9) Enil)) T4 with 
         | Ecall a b c => 
(fun (e0 : expr) (e1 : exprlist) (t0 : type) =>
    get_bit_reg = Ecall e0 e1 t0 ->
    v = Vint (Arm6_State.reg_content s d) [n31]) a b c
 | _ => True end). cbv beta.
  case_I gb_expr. red.
*)

(*
  generalize (refl_equal get_bit_reg).
  pattern get_bit_reg at 1.*)

  (*match goal with [ |- ?concl _ _ _ ] =>
    change 
      (match Ecall a1 a2 a3 with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  
  unfold get_bit_reg in gb_expr.
match goal with [ |- ?concl] => change ((fun _ _ _ => concl) 
   (Evalof (Evar get_bit T16) T16)
   (Econs (reg_id adc_compcert.d)
                    (Econs (Eval (Vint (repr 31)) T9) Enil))
   T4) end.
  match goal with [ gb_expr : context c [Ecall ?a1 ?a2 ?a3] |- ?concl _ _ _ ] =>
    change 
      (match Ecall a1 a2 a3 with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  case_I gb_expr. red.
  intros until rargs. intro ty.
  intros until vres.
  intros rf_exp rargs_exp vf_rval targs_vlst Heqtprf Heqfun Heqtpfun fd_funcall.
  
  match goal with [ |- ?concl _ _ _ ] =>
    change 
      (match get_bit_reg with 
         | Ecall a b c => concl a b c | _ => True end) end. cbv beta.
  

  case_eq get_bit_reg. intro
  case get_bit. intro
  unfold get_bit_reg in get_bit.*)
Admitted.




Lemma same_get_reg :
  forall e m0 m0' vargs m l b s d t m' v,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    proc_state_related m e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m get_rd_bit31 t m' v->
    v = Vint ((Arm6_State.reg_content s d) [n31]).
Proof.
  intros until v. intros av bp psrel dfrel get_bit.
  inv get_bit. 
  (*rename H into get_bit_reg_exp, H0 into get_bit_reg_v.
  inv get_bit_reg_exp.*)
  
  (*unfold get_rd_bit31 in H.
  inv_eval_expr m m'.*)

  inv H.
  inv H4. inv H8. inv H9. inv H5.
  
  (** HERE expand function reg *)



  apply same_reg_d with e m2 t1 m1 a1' l b s d in H4;
    [idtac| exact psrel |exact dfrel].
  rewrite H4 in *. 
  inv H13. inv H5. inv H14.
  inv H0. inv H6. inv H2. inv H4.
  (* by explore local env 'e', we know get_bit isn't in local env*)
  assert (e!get_bit=None).
  inv_alloc_vars e.
    simpl. reflexivity.
  (* esl_evar_global *)
  inv H1;[rewrite H in H5;discriminate|idtac].
    (* pass list of argument values vargs0 to get_bit function *)
    (* first arg (reg_content d) *)
    inv H7. 
    (* from H6, we know v' = (Eval (Vint (Arm6_State.reg_content s d)) T1) *)
    inv H6. 
    (* second arg 31 *)
    inv H13. 
    (* from H6, we know v' = (Eval (Vint (repr 31)) T9) *)
    inv H6.
    (* the rest of arg list is nil *)
    inv H14. 
    (* simpl typeof *)
    simpl in H10, H9.
    (*compcert1.9 improves cast definition 
       (sem_cast v1 t1 t2 = Some v2), proofs are simpler
       than before. *)
    (* cast int32 to uint32 is cast_case_neutral,cast the same value to v1 *)
    inv H9.
    (* cast int32 to uint32 is cast_case_neutral,cast the same value to v0 *)
    inv H10.
    (* find symbol get_bit in global env, return the value of its block b0 *)
    unfold Genv.find_symbol in H4;simpl in H4.
    injection H4;intro;rewrite<-H0 in *;clear H0 H4 H8 b0.
    (* find function in block -7 in global env*)
    rewrite Genv.find_funct_find_funct_ptr in H11.
    unfold Genv.find_funct_ptr in H11. unfold ZMap.get in H11.
    simpl in H11. unfold ZMap.set in H11. simpl in H11. 
    rewrite PMap.gso in H11;[idtac|simpl;congruence].
    unfold PMap.get in H11; simpl in H11.
    injection H11;intro;rewrite<-H0 in *;clear H0 H11 H12 fd.
    (* expand get_bit *)
    (* eval_funcall from m3 to m' *)
    inv H16. 
    (* exec_stmt from m4 to m5 *)
    inv H5.
    simpl in H6.
    (* eval_expression from m4 to m5*)
    inv H10. 
    (* eval Ebinop will split binop with 2 params, m4->m'0;m'0->m5*)
    inv H0.
    (* eval Eval, m4 = m'0*)
    inv H18.
    (* eval Ebinop m4 -> m5,split the two params shr m4->m'0;m'0->m5*)
    inv H17.
    (* eval Evalof, m4 -> m'0*)
    inv H16. 
    (* eval Eval, m4=m'0 *)
    inv H11.
    (* eval Evalof, m'0 -> m5*)
    inv H18. 
    (* eval Evar, m'0=m5 *)
    inv H11.
    (* first param of binop and *)
    (* esr_binop in m5 *)
    inv H5. simpl in H14.
    (* esr_rval in m5, v2 = (Eval (Vint (repr 1)) T9) *)
    inv H13.
    (* second param of binop and *)
    (* esr_binop in m5 *)
    inv H12. simpl in H15.
    (* eval the value of varible x *)
    (* get local env e0 from alloc_variables in m1 *)
    inv_alloc_vars e0.
    (* get the initial value of params x in m5 *)
    inv_bind_params m5. 
    (* the block which contents x, b1 = b2 *)
    injection eget;intro;rewrite<-H0 in *;clear H0 eget b2.
    (* the block which contents n, b0 = b3 *)
    injection eget0;intro;rewrite<-H0 in *;clear H0 eget0 b3.
    (* evaluate the simple expression on value of x *)
    inv H11. 
    (* x is in local env *)
    inv H4;[idtac|simpl in H7;discriminate H7].
    (* block which contents x, b1 = b2*)
    simpl in H11;injection H11;intro;rewrite<-H0 in *;clear H0 H11 H5 b2.
    (* b1 is not changed in m5 and m6 *)    
    unfold store_value_of_type in *; simpl in str, str0.
    unfold load_value_of_type in *; simpl in H9.
    val_not_changed_str AST.Mint32 b1 (0 mod modulus) m6 m5.
    rewrite str0 in H9; clear str0.
    intro str0;generalize str;intro str16.
    eapply Mem.load_store_same in str16;[idtac|simpl;auto].
    (* v2 = (Vint (Arm6_State.reg_content s d))*)
    rewrite str16 in H9;clear str16;simpl in H9.
    injection H9;intro;rewrite<-H0 in *;clear H9 H0 v2.
    (*get the initial value of params n in m5 *)
    (* esr_valof in m5 *)
    inv H13.
    (* esl_var_local in m5, n is in local env *)
    inv H4;[idtac|simpl in H7;discriminate H7].
    (* block which contents n, b1 = b2*)
    simpl in H11;injection H11;intro;rewrite<-H0 in *;clear H0 H11 H5 b2.
    (* load the same value as stored in m6 *)
    unfold load_value_of_type in *; simpl in H9.
    eapply Mem.load_store_same in str0;[idtac|simpl;auto].
    (* v3 = (Vint (repr 31))*)
    rewrite H9 in str0;clear H9.
    injection str0;intro;rewrite H0 in *;clear H0 str0 v3.
    (* calculate v1 the result of sem_shr *)
    unfold sem_shr in H15;simpl in H15.
    injection H15;intro;rewrite<-H0 in *;clear H15 H0 v1.
    (* calculate v0 the result of sem_and *)
    unfold sem_and in H14;simpl in H14.
    injection H14;intro;rewrite<-H0 in *;clear H14 H0 v0.
    (* calculate v the final result *)
    destruct H6. unfold sem_cast in H2;simpl in H2.
    injection H2;intro;rewrite<-H4 in *;clear H2 H4 v.
    (* have hypothesis 0<31<wordsize *)
    assert (wdsz:0<31<Z_of_nat wordsize). unfold wordsize. 
    unfold Wordsize_32.wordsize.
    simpl Z_of_nat. omega.
    rewrite (same_getbit (Arm6_State.reg_content s d) wdsz); reflexivity.
Qed.



Unset Implicit Arguments.
(* Assume that every function that ADC calls, executes correctly
   and the C proc and ARM state related after these function execution *)
Axiom functions_behavior_ok:
  forall e l b s vf fd m vargs t m' vres l' b' s',
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    Genv.find_funct (Genv.globalenv prog_adc) vf = Some fd ->
    eval_funcall (Genv.globalenv prog_adc) m fd vargs t m' vres ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l' b' s')).

(* Assume that call to unpredictable leads to an Ko result*)
Axiom funct_unpredictable:
  forall e semstt vf fd m vargs t m' vres,
    proc_state_related (of_mem proc m) e (Ok tt semstt) ->
    Genv.find_funct (Genv.globalenv prog_adc) vf = Some fd ->
    eval_funcall (Genv.globalenv prog_adc) m fd vargs t m' vres ->
    proc_state_related (of_mem proc m') e 
    (unpredictable Arm6_Message.EmptyMessage semstt).

(* Assume function reg_n only load from memory, not change it*)
Axiom get_reg_ok :
  forall e id m t m' r,
    eval_expr (Genv.globalenv prog_adc) e m RV (reg_id id) t m' r ->
    eval_expr (Genv.globalenv prog_adc) e m RV (reg_id id) t m r/\m=m'.


Definition oldrn_assgnt := 
  Eassign (Evar old_Rn T1) (reg_id n) T1.

(* Assum the assignment of old_Rn has no effect on the part of memory
   where located proc*)
Axiom set_oldrn_ok:
  forall m m' v oldrn_blk ofs,
    store_value_of_type T1 m oldrn_blk ofs v = Some m'->
    of_mem proc m = of_mem proc m'.

Lemma oldrn_assgnt_ok:
 forall e m l b s t m' v,
  proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
  eval_expression (Genv.globalenv prog_adc) e m
    oldrn_assgnt t m' v ->
  proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)).
Proof.
  intros until v. intros psrel rn_as.
  
  inv rn_as. inv H. inv H4.
  eapply get_reg_ok in H5. inv H5.
  simpl in *.
  eapply set_oldrn_ok in H11.
  
  rewrite <- H11. exact psrel.
Qed.

(* Lemmas on if ConditionPassed*)
Definition condpass :=
  Ecall (Evalof (Evar ConditionPassed T5) T5)
  (Econs
    (Eaddrof
      (Efield (Ederef (Evalof (Evar proc T3) T3) T6) cpsr
        T7) T8) (Econs (Evalof (Evar cond T9) T9) Enil))
  T10.

Axiom no_effect_condpass :
  forall e m m' t v,
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->    
    m = m'.


(* try with external function ConditionPassed, failed *)
(*Lemma condpass_bool' :
  forall m0 m0' m0'' vargs e bcond m t m' v cd l bo s b,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->    
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m0'' ->
    e!cond=Some (bcond,Tint I32 Signed) ->
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->
    Mem.load AST.Mint32 m0'' bcond (0 mod modulus) = 
    Mem.load AST.Mint32 m bcond (0 mod modulus)->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l bo s)) ->
    cond_func_related m' e cd ->
    bool_val v T4 = Some b ->
    Arm6_Functions.State.ConditionPassed s cd = b.
Proof.
  intros.
  unfold cond_func_related in H5. unfold cond_proj in H5.
  unfold varg_proj in H5. unfold param_val in H5.
  (* alloc_variables gives the info on variable allocation on blocks *)
  Set Printing Depth 50.
  
  generalize H1;intro econd. 
  inv_alloc_vars e. simpl. 
  simpl in H1;injection H1;intro;subst;clear H1.
  pose (e:= (PTree.set old_Rn (b6, Tint I32 Unsigned)
            (PTree.set shifter_operand (b5, Tint I32 Unsigned)
               (PTree.set n (b4, Tint I8 Unsigned)
                  (PTree.set d (b3, Tint I8 Unsigned)
                     (PTree.set cond (bcond, Tint I32 Signed)
                        (PTree.set S (b0, Tint I8 Signed)
                           (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                              empty_env))))))));
  fold e in H0, H2, H4, econd.
  (* bind_parameters gives the info on initial value of parameters and storage 
     block *)
  inv_bind_params m0''.
  injection eget; intro; rewrite<-H in *;clear H eget b2;
  injection eget0; intro; rewrite<- H in *;clear H eget0 b7;
  injection eget1; intro; rewrite<- H in *;clear H eget1 b8;
  injection eget2; intro; rewrite<- H in *;clear H eget2 b9;
  injection eget3; intro; rewrite<- H in *;clear H eget3 b10;
  injection eget4; intro; rewrite<- H in *;clear H eget4 b11.

  unfold store_value_of_type in *;
  simpl in str, str0, str1, str2, str3, str4.

  (*value in b2 is not changed between m10 and m0'' *)
  val_not_changed_str AST.Mint32 bcond (0 mod modulus) m10 m0''.
  intros str5 str6 str7.
  rewrite str2 in str3; clear str2.
  rewrite str3 in str4; clear str3.
  (* load_store the same for the value of b2 in m10 *)
  apply Mem.load_store_same in str1;[idtac|admit(*TODO*)].
  rewrite H3 in str4; clear H3.
  rewrite<-str4 in str1; clear str4.
  unfold load_value_of_type;simpl.
  (* from eval_expression condpass , m = m' *)
  apply no_effect_condpass in H2.
  destruct H2.
  rewrite H in *;clear H m.
  (* relation between v and b *)
  rewrite str1. simpl.
  (* in C, the relation between v2 and v, how to calculate v from v2 *)
  (* eval_expression -> eval_expr, from m to m' *)
  inv H0.
  (* eval_funcall, from m to m' *)
  inv H.
  (* eval_evalof, from m' to m1 *)
  inv H5.
  (* eval_evar, m' = m1 *)
  inv H11.
(* in new version of CompCert1.9, there are several changes in semantic definition
   which have influence on our proof.*)
  (* v = vres *)
  inv H1.
  (* esr_valof in m13 *)
  inv H8. 
  (* esl_val_global *)
  inv H1;[discriminate|idtac].
  (* find ConditionPassed in global *)
  unfold Genv.find_symbol in H8;  simpl in H8.
  injection H8;intro;rewrite<-H in *;clear H8 H b2 H3.
  unfold load_value_of_type in H5;simpl in H5.
  injection H5;intro;rewrite<-H in *;clear H5 H vf.
  simpl in H13. 
  destruct eq_dec;[idtac|discriminate].
  (* clear useless Hyp *)
  clear e0 H2 H15 H14.
  (* fd is the external function ConditionPassed *)
  inversion H13;clear H13. rewrite<-H0 in *;clear H0.
  (* pass params to ConditionPassed *)
  (* first param proc->cpsr *)
  inv H7.
  (* eval_addrof, from m1 to m14 *)
  inv H3. 
  (* eval_field, from m1 to m14 *)
  inv H5. 
  (* eval_deref, from m1 to m14 *)
  inv H13. 
  (* eval_valof, from m1 to m14 *)
  inv H3. 
  (* eval_var, m1=m14 *)
  inv H5.
  (* second param cond *)
  inv H12.
  (* eval_valof, from m14 to m1 *)
  inv H3.
  (* eval_var, m14=m1 *)
  inv H5.
  (* no more params *)
  inv H11.
  (* value of first param proc->cpsr *)
  inv H9. simpl in H2. simpl in H10.
  injection H10;intros; subst;clear H10.
  (* esr_addrof in m13 *)
  inv H1.
  unfold sem_cast in H2;simpl in H2.
  injection H2;intro;subst;clear H2.
  (* value of first param is Vptr b2 ofs *)
  (* get the value of b2 and ofs in m13 *)
  (* esl_field_struct in m13*)
  inv H5;[idtac|discriminate].
  injection H9;intros Hid0 Hfl;rewrite<-Hfl in *;rewrite<-Hid0 in *;
  clear H9 Hid0 Hfl.
  apply field_offset_in_range 
    with SLv6_Processor _ _ _ typ_SLv6_StatusRegister in H10;
  [idtac|simpl;
  repeat(destruct AST.ident_eq;discriminate||(try reflexivity)
    ||(try (destruct n0;reflexivity)))].
  (* esl_deref in m12 *)
  inv H2.
  (* esr_rvalof in m12 *)
  inv H5.
  (* esl_var_local in m12 *)
  inv H1;[simpl in H9;injection H9;intros Hp;rewrite<-Hp in *;clear b7 Hp H9 H2
    |simpl in H3;discriminate].
  (* value of second param cond *)
  inv H7. simpl in H9.
  (* esr_valof in m12 *)
  inv H3. clear H2.
  (* find cond in local env *)
  (* esl_var_local in m14 *)
  inv H1;[rewrite econd in H5;injection H5;intro;rewrite<-H in *;clear econd H H5 b7
    |rewrite econd in *;discriminate].
  (* v'= Val.load_result AST.Mint32 v2*)
  unfold load_value_of_type in H7;simpl in H7;
  rewrite str1 in H7;clear str1.
  injection H7;intro Hv;rewrite<-Hv in *;clear Hv H7.
  unfold sem_cast in H9;simpl in H9.
  (* no more param *)
  inv H11.
  (* eval_funcall, from m13 to m13 *)
  inv H18.
  (* external_call from m13 to m13 *)
  inv H12.
  (* first event value *)
  inv H.
  (* second event value *)
  inv H13.
  (* no more event *)
  inv H14.
  (* Translation between values and event values. *)
  (* v6 can be either a Vint or a Vptr *)
  destruct v2;[discriminate
    |injection H9;intro Hi;rewrite<-Hi in *;clear H9 Hi v6
    |discriminate
    |injection H9;intro Hb;rewrite<-Hb in *;clear H9 Hb v6].
    (* v2 is Vint *)
    inv H0.
*)

Lemma condpass_bool :
  forall m0 m0' e m t m' v cond s b,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    eval_expression (Genv.globalenv prog_adc) e m condpass t m' v ->
    bool_val v T4 = Some b ->
    Arm6_Functions.State.ConditionPassed s cond = b.
Proof.
Admitted.

(*Lemma on proc_state_relates holds after set_reg*)
Definition set_regpc :=
  Ecall (Evalof (Evar set_reg_or_pc T11) T11)
  (Econs (Evalof (Evar proc T3) T3)
    (Econs (Evalof (Evar d T4) T4)
      (Econs
        (Ebinop Oadd
          (Ebinop Oadd
            (Evalof (Evar old_Rn T1) T1)
            (Evalof (Evar shifter_operand T1) T1)
            T1)
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T10) T10)
          T10) Enil))) T12.

Lemma same_setregpc :
  forall e m l b s0 s t m' v d n so ,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    eval_expression (Genv.globalenv prog_adc) e m set_regpc t m' v ->
    (forall l b, proc_state_related (of_mem proc m') e 
      (Ok tt (mk_semstate l b
        (Arm6_State.set_reg s d (add (add (Arm6_State.reg_content s0 n) so)
          ((Arm6_State.cpsr s)[Cbit]) ))))).
Proof.
  intros until so. intros psrel setreg. intros.
  inv setreg. inv H. inv H4. inv H9. inv H5. inv H4. inv H5.
  inv H14. inv H4. inv H5. inv H13. inv H4. inv H17. inv H15. inv H4.
  inv H19. inv H4. inv H18. inv H4. inv H15. inv H13. inv H4. inv H5.
  inv H14. inv H0.
Admitted.


(* Lemmas on if S==1 *)

Definition is_S_set :=
  Ebinop Oeq (Evalof (Evar S T10) T10)
    (Eval (Vint (repr 1)) T9) T9.

Lemma no_effect_is_S_set :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v ->
    m = m'.
Proof.
  intros until v. intros is_s. 
  inv is_s. unfold is_S_set in H.  
  inv_eval_expr m m'.
  reflexivity.
Qed.

Lemma S_bool :
  forall m0 e m0' m t m' v sbit b,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    sbit_func_related m e sbit ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set t m' v ->
    bool_val v T9 = Some b->
    Util.zeq sbit 1 = b.
Proof.
  intros until b. intros av sfrel ee bv.
  unfold sbit_func_related in sfrel. unfold bit_proj in sfrel.
  unfold param_val in sfrel.
  inv_alloc_vars e;
  pose (e:=
    (PTree.set old_Rn (b6, Tint I32 Unsigned)
      (PTree.set shifter_operand (b5, Tint I32 Unsigned)
        (PTree.set n (b4, Tint I8 Unsigned)
          (PTree.set d (b3, Tint I8 Unsigned)
            (PTree.set cond (b2, Tint I32 Signed)
              (PTree.set S (b0, Tint I8 Signed)
                (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                  empty_env))))))));
  fold e in ee;simpl.
  (* eval_expression is_S_set from m to m' *)
  inv ee. unfold is_S_set in H.
  (* eval_expr from m to m' *)
  inv_eval_expr m m'.
  (* params of binop eq *)
  (* esr_binop in m' *)
  inv esr. simpl in H6.
  (* S *)
  (* esr_valof in m' *)
  inv H4. clear H2.
  (* esl_var_local in m' *)
  inv H1;[simpl in H4;injection H4;intro Heq;rewrite<-Heq in *;clear b7 Heq H4
    |discriminate].
  (* v6 is the value of S in m' *)
  unfold T10 in H7;simpl in H7;rewrite H7.
  (* esr_rval in m' *)
  inv H5.
  (* v1 is either Vint of Vptr *)
  destruct v1;
    [discriminate
      |unfold sem_cmp in H6;simpl in H6;
        injection H6;intro Heq;rewrite<-Heq in *;clear Heq H6 v
      |discriminate
      |discriminate].
  unfold varg_proj.
  unfold bool_val in bv;simpl in bv.
  unfold w1.
  destruct (eq i (repr 1));
  simpl in bv;injection bv;intro;rewrite<-H;clear H bv b;
  reflexivity.
Qed.

(* Lemmas on if (((S == 1) && (d == 15)))*)
Definition is_S_set_and_is_pc :=
  Econdition
  (Ebinop Oeq (Evalof (Evar S T10) T10)
    (Eval (Vint (repr 1)) T9) T9)
  (Econdition
    (Ebinop Oeq (Evalof (Evar d T4) T4)
      (Eval (Vint (repr 15)) T9) T9)
    (Eval (Vint (repr 1)) T9)
    (Eval (Vint (repr 0)) T9) T9)
  (Eval (Vint (repr 0)) T9) T9.


Lemma no_effect_is_S_set_and_is_pc :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v ->
    m = m'.
Proof.
  intros until v. intro ee.
  inv ee.
  unfold is_S_set_and_is_pc in H.
  inv_eval_expr m m'.
  destruct b.
    (*b1 true*)
    inv_eval_expr m'0 m'.
    destruct b.
      (*b2 true*)
      inv_eval_expr m'1 m'.
      reflexivity.
      (*b2 false*)
      inv_eval_expr m'1 m'.
      reflexivity.
    (*b1 false*)
    inv_eval_expr m'0 m'.
    reflexivity.
Qed.

Lemma same_reg_val :
forall x y,
  (eq x (repr y) = Util.zeq (mk_regnum x) y).
Proof.
Admitted.

Lemma S_pc_bool :
  forall e m t m' v sbit d b,
    sbit_func_related m e sbit ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m is_S_set_and_is_pc t m' v ->
    bool_val v T9 = Some b ->
    Util.zeq sbit 1 && Util.zeq d 15 = b.
Proof.
Admitted.

(*Ltac inv_eval_simple m ex :=
  match goal with
    |[eslst:eval_simple_list ?ge ?e m (Econs ?r ?rl) ?tylst ?vlst|-?cl]=>
      inv eslst;inv_eval_simple m r;inv_eval_simple m rl
    |[eslst:eval_simple_list ?ge ?e m Enil ?t ?rl|-?cl]=>
      inv eslst
    |[esl:eval_simple_lvalue ?ge ?e m (Eloc ?b1 ?ofs1 ?ty) ?b2 ?ofs2|-?cl]=>
      inv esl
    |[esl:eval_simple_lvalue ?ge ?e m (Evar ?x ?ty) ?b ?ofs|-?cl]=>
      inv esl;[try discriminate|try discriminate]
    |[esl:eval_simple_lvalue ?ge ?e m (Ederef ?r ?ty) ?b ?ofs|-?cl]=>
      inv esl;inv_eval_simple r m
    |[esl:eval_simple_lvalue ?ge ?e m (Efield ?l ?f ?ty) ?b ?ofs|-?cl]=>
      inv esl;inv_eval_simple l m
    |[esr:eval_simple_rvalue ?ge ?e m (Eval ?vres ?ty) ?v|-?cl]=>
      inv esr
    |[esr:eval_simple_rvalue ?ge ?e m (Evalof ?l ?ty) ?v|-?cl]=>
      inv esr;inv_eval_simple m l
    |[esr:eval_simple_rvalue ?ge ?e m (Eaddrof ?l ?ty) ?v|-?cl]=>
      inv esr;inv_eval_simple m l
    |[esr:eval_simple_rvalue ?ge ?e m (Eunop ?op ?r1 ?ty) ?v|-?cl]=>
      inv esr;inv_eval_simple m r1
    |[esr:eval_simple_rvalue ?ge ?e m (Ebinop ?op ?r1 ?r2 ?ty) ?v|-?cl]=>
      inv esr;inv_eval_simple m r1;inv_eval_simple m r2
    |[esr:eval_simple_rvalue ?ge ?e m (Ecast ?r1 ?ty) ?v|-?cl]=>
      inv esr;inv_eval_simple m r1
    |[esr:eval_simple_rvalue ?ge ?e m (Esizeof ?ty1 ?ty) ?v|-?cl]=>
      inv esr
  end.
*)
Ltac inv_eval_simple m ex :=
  match goal with
    |[eslst:eval_simple_list ?ge ?e m ex ?tylst ?vlst|-?cl]=>
      match ex with
        |Econs ?r ?rl=>inv eslst;inv_eval_simple m r;inv_eval_simple m rl
        |Enil=>inv eslst
      end
    |[esl:eval_simple_lvalue ?ge ?e m ex ?b ?ofs|-?cl]=>
      match ex with
        |Eloc ?b1 ?ofs1 ?ty=>inv esl
        |Evar ?x ?ty=>inv esl;[try discriminate|try discriminate]
        |Ederef ?r ?ty=>inv esl;inv_eval_simple m r
        |Efield ?l ?f ?ty=>inv esl;inv_eval_simple m l
      end
    |[esr:eval_simple_rvalue ?ge ?e m ex ?v|-?cl]=>
      match ex with
        |Eval ?vres ?ty=>inv esr
        |Evalof ?l ?ty=>inv esr;inv_eval_simple m l
        |Eaddrof ?l ?ty=>inv esr;inv_eval_simple m l
        |Eunop ?op ?r1 ?ty=>inv esr;inv_eval_simple m r1
        |Ebinop ?op ?r1 ?r2 ?ty=>
          inv esr;inv_eval_simple m r1;inv_eval_simple m r2
        |Ecast ?r1 ?ty=>inv esr;inv_eval_simple m r1
        |Esizeof ?ty1 ?ty=>inv esr
      end
  end.


(* Lemmas on if CurrentModeHasSPSR *)
Definition hasSPSR :=
  Ecall (Evalof (Evar CurrentModeHasSPSR T13) T13)
  (Econs (Evalof (Evar proc T3) T3) Enil) T10.


Lemma if_hasSPSR_ok' :
  forall m0 e m0' m t m' v id ty,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    Mem.nextblock m0' < Mem.nextblock m ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    In (id,ty) (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars))->
    param_val id m e=param_val id m' e.
Proof.
  intros until ty. intros av mn ee inlst.
  inv ee. unfold hasSPSR in H.
  (* eval_expr between m and m' *)

  inv_eval_expr m m'.

  (* alloc_vars *)
  inv_alloc_vars e.
  pose (e:=(PTree.set old_Rn (b6, Tint I32 Unsigned)
            (PTree.set shifter_operand (b5, Tint I32 Unsigned)
               (PTree.set n (b4, Tint I8 Unsigned)
                  (PTree.set d (b3, Tint I8 Unsigned)
                     (PTree.set cond (b2, Tint I32 Signed)
                        (PTree.set S (b0, Tint I8 Signed)
                           (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                              empty_env))))))));
  fold e in esr0, esr1, esr; fold e.
  (* esr in m', v is vres *)
  inv_eval_simple m' (Eval vres T10).
  (* esr in m3, find vf is CurrentModeHasSPSR *)
  inv_eval_simple m2 ((Evalof (Evar CurrentModeHasSPSR T13) T13)).
  (* find block b *)
  unfold Genv.find_symbol in H5;simpl in H5.
  injection H5;intro;rewrite<-H in *;clear H b H5 H8 H2.
  unfold load_value_of_type in H4;simpl in H4;
    injection H4;intro;rewrite<-H in *;clear H vf H4.
  (* fd is in block -6, and it is CurrentModeHasSPSR *)
  rewrite Genv.find_funct_find_funct_ptr in Heqff.
  unfold Genv.find_funct_ptr in Heqff;unfold ZMap.get in Heqff;simpl in Heqff.
  unfold ZMap.set in Heqff;simpl in Heqff. 
  repeat (rewrite PMap.gso in Heqff;[idtac|simpl;congruence]).
  rewrite PMap.gss in Heqff.
  injection Heqff;intro;rewrite<-H in *;clear H Heqff fd.
  (* pass variable proc to eval_function *)
  inv_eval_simple m2 (Econs (Evalof (Evar proc T3) T3) Enil).
  (* type of ty*)
  injection Heqtf;intros Htres Hty;rewrite<-Htres in *;rewrite<-Hty in *;
    clear Heqtf Hty Htres ty0 tres H5 Heqcf.
  (* cast v' into v0 *)
  simpl in H2;unfold sem_cast in H2;simpl in H2.
  (* eval_funcall from m3 to m' *)
  inv ev_funcall.
  (* exec_stmt from m9 to m10 *)
  inv H5. simpl in H6.
  (* eval_expression from m9 to m10 *)
  inv H12.
  (* eval_expr from m9 t m10 *)
  inv_eval_expr m9 m10.
  (* free_list from m10 to m' *)
  inv_alloc_vars e0.
  simpl in alc6, alc5.
  (* Mem.free from m10 to m'*)
  assert(Mem.free m10 b7 0 4 = Some m').
  simpl in H10;rewrite<-H10;
  destruct (Mem.free m10 b7 0 4); reflexivity.
  (* the parameter list *)
  unfold In in inlst;simpl in inlst.
  (*b=b1*)
  simpl in H9;injection H9;intro eq;rewrite<-eq in *;clear H9 eq b.
  (* b6<b7 *)
  generalize alc6 alc5;intros alc6' alc5'.
  apply Mem.alloc_result in alc6';
  apply Mem.valid_new_block in alc5';
  unfold Mem.valid_block in alc5';
  rewrite<-alc6' in mn;
  apply (Zlt_trans b6) in mn;[idtac|exact alc5'];
  clear alc6' alc5'.

  (* case on parameters *)
  destruct inlst as [param|[param|[param|[param|[param|[param|[param|inlst]]]]]]];
  try
  (injection param;intros Hptp Hpid;rewrite<-Hpid;clear Hptp Hpid param id0 ty;
  (* simplify in goal *)
  unfold param_val;simpl;
  unfold load_value_of_type in *;simpl in H8 |-*);
  (* bind parameters from m8 to m10 *)
  inv_bind_params m10; repeat rrw_block;
  unfold store_value_of_type in str;simpl in str.

  (* param proc *)
  (* load b1 from m2 is v' *)
  rewrite H8.
  
  (* stores between m8 and m10 do not change value in b1 *)
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint32 b1 (0 mod modulus) in str;
    [idtac|left;blocks_lt b1 b6;blocks_neq b1 b7;exact mn].
  (* load the same value in b1 from m10 to m' *)
  rewrite Mem.load_free with m10 b7 0 4 m' AST.Mint32 b1 (0 mod modulus);
    [idtac|exact H|left;blocks_lt b1 b6;blocks_neq b1 b7;exact mn].
  (* load same value in b1 from m2 and m8*)
  rewrite Mem.load_alloc_other with
    m2 0 4 m8 b7 AST.Mint32 b1 (0 mod modulus) v' in str;
    [rewrite str;reflexivity|exact alc6|exact H8].
  (*
  (* b1<>b7*)
  assert(Hneqb17:b1<>b7).
  (* b1<b6 *)
  blocks_lt b1 b6.
  (* b1 <> b7*)
  blocks_neq b1 b7.
  exact mn.
  (* load the same value in b1 from m10 to m' *)
  assert
    (ld10':Mem.load AST.Mint32 m' b1 (0 mod modulus)
      =Mem.load AST.Mint32 m10 b1 (0 mod modulus)).
  apply Mem.load_free with b7 0 4;
    [exact H|left;exact Hneqb17].
  (* stores between m8 and m10 do not change value in b1 *)
  inv_bind_params m10; repeat rrw_block.
  unfold store_value_of_type in str;simpl in str.
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint32 b1 (0 mod modulus) in str;
  [idtac|left;exact Hneqb17].
  rewrite str in ld10';clear str.
  (* load same value in b1 from m3 and m8*)
  simpl in alc6;
  apply Mem.load_alloc_other with 
    m2 0 4 m8 b7 AST.Mint32 b1 (0 mod modulus) v' in alc6;[idtac|exact H8].
  (* load same value in b1 from m8 to m' *)
  rewrite alc6 in ld10';clear alc6.
  rewrite ld10';reflexivity.*)

  (* param S *)
  (* stores between m8 and m10 do not change value in b0 *)
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint8signed b0 (0 mod modulus) 
    in str;
    [idtac|left;blocks_lt b0 b6;blocks_neq b0 b7;exact mn].
  (* load the same value in b0 from m10 to m' *)
  rewrite Mem.load_free with m10 b7 0 4 m' AST.Mint8signed b0 (0 mod modulus);
    [idtac|exact H|left;blocks_lt b0 b6;blocks_neq b0 b7;exact mn].
  (* load same value in b0 from m2 and m8*)
  rewrite Mem.load_alloc_unchanged with
    m2 0 4 m8 b7 AST.Mint8signed b0 (0 mod modulus) in str;
    [rewrite str;reflexivity|exact alc6
      |unfold Mem.valid_block;apply Mem.alloc_result in alc6;
        rewrite<-alc6;blocks_lt b0 b6;blocks_lt' b0 b7;exact mn].
  (*
  (* b0<b7*)
  assert(Hltb07:b0<b7).
  blocks_lt b0 b6;blocks_lt' b0 b7. exact mn.
  generalize Hltb07;intro Hneqb07;apply Zlt_not_eq in Hneqb07.
  (* load the same value in b0 from m10 to m' *)
  assert
    (ld10':Mem.load AST.Mint8signed m' b0 (0 mod modulus)
      =Mem.load AST.Mint8signed m10 b0 (0 mod modulus)).
  apply Mem.load_free with b7 0 4;
    [exact H|left;exact Hneqb07].
  (* stores between m8 and m10 do not change value in b0 *)
  inv_bind_params m10; repeat rrw_block.
  unfold store_value_of_type in str;simpl in str.
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint8signed b0 (0 mod modulus) 
    in str;
  [idtac|left;exact Hneqb07].
  rewrite str in ld10';clear str.
  (* load same value in b0 from m3 and m8*)
  simpl in alc6;
  apply Mem.load_alloc_unchanged with 
    m2 0 4 m8 b7 AST.Mint8signed b0 (0 mod modulus) in alc6;
    [rewrite alc6 in ld10';clear alc6;rewrite ld10';reflexivity
      |unfold Mem.valid_block;apply Mem.alloc_result in alc6;
        rewrite<-alc6;exact Hltb07].*)

  (* param cond *)
  (* stores between m8 and m10 do not change value in b2 *)
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint32 b2 (0 mod modulus) 
    in str;
    [idtac|left;blocks_lt b2 b6;blocks_neq b2 b7;exact mn].
  (* load the same value in b2 from m10 to m' *)
  rewrite Mem.load_free with m10 b7 0 4 m' AST.Mint32 b2 (0 mod modulus);
    [idtac|exact H|left;blocks_lt b2 b6;blocks_neq b2 b7;exact mn].
  (* load same value in b2 from m2 and m8*)
  rewrite Mem.load_alloc_unchanged with
    m2 0 4 m8 b7 AST.Mint32 b2 (0 mod modulus) in str;
    [rewrite str;reflexivity|exact alc6
      |unfold Mem.valid_block;apply Mem.alloc_result in alc6;
        rewrite<-alc6;blocks_lt b2 b6;blocks_lt' b2 b7;exact mn].
  (*
  (* b2<b7*)
  assert(Hltb27:b2<b7).
  blocks_lt b2 b6;blocks_lt' b2 b7;exact mn.
  generalize Hltb27;intro Hneqb27;apply Zlt_not_eq in Hneqb27.
  (* load the same value in b2 from m10 to m' *)
  assert
    (ld10':Mem.load AST.Mint32 m' b2 (0 mod modulus)
      =Mem.load AST.Mint32 m10 b2 (0 mod modulus)).
  apply Mem.load_free with b7 0 4;[exact H|left;exact Hneqb27].
  (* stores between m8 and m10 do not change value in b2 *)
  inv_bind_params m10; repeat rrw_block.
  unfold store_value_of_type in str;simpl in str.
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint32 b2 (0 mod modulus) 
    in str;
  [idtac|left;exact Hneqb27].
  rewrite str in ld10';clear str.
  (* load same value in b0 from m3 and m8*)
  simpl in alc6;
  apply Mem.load_alloc_unchanged with 
    m2 0 4 m8 b7 AST.Mint32 b2 (0 mod modulus) in alc6;
    [rewrite alc6 in ld10';clear alc6;rewrite ld10';reflexivity
      |unfold Mem.valid_block;apply Mem.alloc_result in alc6;
        rewrite<-alc6;exact Hltb27].*)
  
  (* parameter d *)
  admit.
  (* parameter n *)
  admit.
  (* parameter shifter_operand *)
  admit.
  (* local variable old_Rn *)
  admit.
  (* parameter list is nil *)
  contradiction.
Qed.

Lemma if_hasSPSR_ok'' :
  forall m0 e m0' m t m' v,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    Mem.nextblock m0' < Mem.nextblock m ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    (exists i, param_val i m e=param_val i m' e).
Proof.
  intros until v. intros av mn ee.
  inv ee. unfold hasSPSR in H.
  (* eval_expr between m and m' *)
  inv_eval_expr m m'.
  (* alloc_vars *)
  inv_alloc_vars e.
  pose (e:=(PTree.set old_Rn (b6, Tint I32 Unsigned)
            (PTree.set shifter_operand (b5, Tint I32 Unsigned)
               (PTree.set n (b4, Tint I8 Unsigned)
                  (PTree.set d (b3, Tint I8 Unsigned)
                     (PTree.set cond (b2, Tint I32 Signed)
                        (PTree.set S (b0, Tint I8 Signed)
                           (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                              empty_env))))))));
  fold e in esr0, esr1, esr; fold e.
  (* esr in m', v is vres *)
  inv_eval_simple m' (Eval vres T10).
  (* esr in m3, find vf is CurrentModeHasSPSR *)
  inv_eval_simple m2 ((Evalof (Evar CurrentModeHasSPSR T13) T13)).
  (* find block b *)
  unfold Genv.find_symbol in H5;simpl in H5.
  injection H5;intro;rewrite<-H in *;clear H b H5 H8 H2.
  unfold load_value_of_type in H4;simpl in H4;
    injection H4;intro;rewrite<-H in *;clear H vf H4.
  (* fd is in block -6, and it is CurrentModeHasSPSR *)
  rewrite Genv.find_funct_find_funct_ptr in Heqff.
  unfold Genv.find_funct_ptr in Heqff;unfold ZMap.get in Heqff;simpl in Heqff.
  unfold ZMap.set in Heqff;simpl in Heqff.
  repeat (rewrite PMap.gso in Heqff;[idtac|simpl;congruence]).
  rewrite PMap.gss in Heqff.
  injection Heqff;intro;rewrite<-H in *;clear H Heqff fd.
  (* pass variable proc to eval_function *)
  inv_eval_simple m2 (Econs (Evalof (Evar proc T3) T3) Enil).
  (* type of ty*)
  injection Heqtf;intros Htres Hty;rewrite<-Htres in *;rewrite<-Hty in *;
    clear Heqtf Hty Htres ty tres Heqcf.
  (* cast v' into v0 *)
  simpl in H2;unfold sem_cast in H2;simpl in H2.
  (* eval_funcall from m3 to m' *)
  inv ev_funcall.
  (* exec_stmt from m9 to m10 *)
  inv H6. simpl in H7.
  (* eval_expression from m9 to m10 *)
  inv H13.
  (* eval_expr from m9 t m10 *)
  inv_eval_expr m9 m10.
  (* free_list from m10 to m' *)
  inv_alloc_vars e0.
  (* Mem.free from m10 to m'*)
  assert(Mem.free m10 b7 0 4 = Some m').
  simpl in H11;rewrite<-H11;
  destruct (Mem.free m10 b7 0 4); reflexivity.
  (* example proc *)
  exists proc.
  (* simplify in goal *)
  unfold param_val. rewrite H9.
  unfold load_value_of_type in *;simpl in H8 |-*.
  rewrite H8.
  (* bind parameters *)
  inv_bind_params m10;rrw_block.
  unfold store_value_of_type in str;simpl in str.
  (* b = b1 *)
  simpl in H9;injection H9;intro Heq;rewrite<-Heq in *;clear H9 Heq b.
  (* b1<>b7*)
  assert(Hneqb17:b1<>b7).
  (* b1<b6 *)
  blocks_lt b1 b6.
  (* b6<b7 *)
  apply Mem.alloc_result in alc6;
  apply Mem.valid_new_block in alc5;
  unfold Mem.valid_block in alc5;
  rewrite<-alc6 in mn.
  apply (Zlt_trans b6) in mn;[idtac|exact alc5].
  (* b1 <> b7*)
  blocks_neq b1 b7.
  exact mn.
  (* stores between m8 and m10 do not change value in b1 *)
  apply Mem.load_store_other with 
    AST.Mint32 m8 b7 (0 mod modulus) v0 m10 AST.Mint32 b1 (0 mod modulus) in str;
    [idtac|left;exact Hneqb17].
  (* load the same value in b1 from m10 to m' *)
  rewrite Mem.load_free with m10 b7 0 4 m' AST.Mint32 b1 (0 mod modulus);
    [idtac|exact H|left;exact Hneqb17].
  (* load same value in b1 from m2 and m8*)
  rewrite Mem.load_alloc_other with
    m2 0 4 m8 b7 AST.Mint32 b1 (0 mod modulus) v' in str;
    [rewrite str;reflexivity|exact alc6|exact H8].
Qed.

Lemma if_hasSPSR_ok :
  forall e m t m' v,
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    m = m'.
Proof.
Admitted.
  

Lemma hasSPSR_true' :
  forall m0 m0' e m vargs t m' v l b s,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)) ->
    bool_val v T4 = Some true ->
    word_of_proc_mode (mode_proj m' e) < 5.
Proof.
Admitted.

(*Lemma hasSPSR_true' :
  forall m0 m0' e m vargs t m' v l b s,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)) ->
    Csem.is_true v T4 ->
    word_of_proc_mode (mode_proj m' e) < 5.
Proof.
  intros until s. intros av bp hs psrel tr.

  inv hs. inv H. inv H0. 
  (* m = m3 *)
  inv H4. inv H3. inv H5. inv H3. inv H4. inv H13.
  (* ? *)
  inv H6.
  (* expand local env e *)
  inv av. inv H14. inv H17. inv H18. inv H19. inv H20. inv H21. inv H22.
  pose (e:=
    PTree.set old_Rn (b7, Tint I32 Unsigned)
      (PTree.set shifter_operand (b6, Tint I32 Unsigned)
        (PTree.set n (b5, Tint I8 Unsigned)
          (PTree.set d (b4, Tint I8 Unsigned)
            (PTree.set cond (b3, Tint I32 Signed)
              (PTree.set S (b2, Tint I8 Unsigned)
                (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                  empty_env))))))).
  fold e in psrel, bp, H7. fold e. 
  (* CurrentModeHasSPSR is in global env *)
  inv H1; [simpl in H6; discriminate H6| clear H3].
  (* search CurrentModeHasSPSR in global env *)
  (* vf=Vptr (-6) w0 *)
  inv H5. unfold load_value_of_type in H4; simpl in H4. 
  injection H4; intro; clear H4. rewrite <- H in *; clear vf H.
  (* fd = fun_Internal_CurrentModeHasSPSR *)
  inversion H11;  destruct eq_dec; 
    [clear e0 H11 H2 H12 H8; inv H0|discriminate H0].

  (* pass parameter proc to internal function CurrentModeHasSPSR *)
  inv H7. inv H5. 
  (* v0 is value of proc *)
  inv H1; clear H4.
  inv H3;
  [unfold e in H5;simpl in H5;injection H5;intro;rewrite<-H in *;clear b0 H H5
  |unfold e in H1;simpl in H1;discriminate H1].


  (* open CrrentModeHasSPSR *)
  inv H16. inv H4. 
  (* return value is v (cast from v1) *)
  simpl in H5; destruct H5.
  (* m9 = m10 *)
  inv H11. inv H5. inv H27. inv H26. inv H16. inv H25. inv H24. inv H16. inv H21.
  (* arguments v2,v3 of binary operation lt*)
  inv H7. simpl in H23.
  (* v3 = 5 *)
  inv H22.
  (* v2 = v0 *)
  inv H21; clear H11.
  (* typ_struct_SLv6_StatusRegister is a structure *)
  inv H9;[idtac|simpl in H24;unfold T7 in H24;discriminate H24].
  inv H24.
  (* offset of mode is 16 *)
  assert (field_offset mode typ_struct_SLv6_StatusRegister = OK 16).  
  unfold field_offset. simpl. 
  Ltac unfold_identeq :=
    destruct AST.ident_eq;
      [try (unfold align;simpl;discriminate||destruct AST.ident_eq)
        |try unfold_identeq].
  unfold_identeq. unfold align. simpl. reflexivity. admit.
  rewrite H5 in H25; clear H5. 
  injection H25;intro;rewrite<-H5 in H16;clear H5 H25 delta.
  (* typ_struct_SLv6_Processor is a structure *)    
  inv H12; [idtac|simpl in H24;unfold T6 in H24;discriminate H24].
  inv H24.
  (* offset of cpsr  is 2 *)
  assert (field_offset cpsr typ_struct_SLv6_Processor = OK 2). admit.
  rewrite H5 in H25; clear H5. 
  injection H25; intro; rewrite<-H5 in H16; clear delta H5 H25.
  (* expand e0 *)
  inv H1. inv H26.   
  (* proc is in e0 *)
  inv H11. inv H12. inv H7;[idtac|simpl in H11; discriminate H11]. clear H9.
  (* b9 = b8 *)
  simpl in H22; injection H22;intro;rewrite<-H1 in *; clear b9 H22 H1.
  (* load v0 from b9 *)
  inv H3.
  inv H28; simpl in H26;injection H26;intro;rewrite<-H1 in *;clear b9 H1 H26.
  unfold store_value_of_type in H27;simpl in H27.
  generalize H27; intro bp'.
  apply Mem.load_store_same in H27;
    [idtac|simpl;destruct v0;simpl;try(exact I||inv H2)].
  unfold load_value_of_type in *; simpl in H6, H16, H21.
  rewrite H27 in H21. 
  injection H21; intro. destruct v0; try discriminate H1.
  injection H1; intros; rewrite<-H3,H5 in *;clear H1 H3 H5.
  simpl in H27.
  (* v' = Vptr b0 i*)
  inv H2.
  unfold sem_cmp in H23; simpl in H23.
  destruct v2; try discriminate H23.
  injection H23; intro; clear H23. rewrite <- H1 in *; clear H1.

  (* unfold goal *)
  unfold mode_proj. unfold find_mode. unfold find_cpsr. unfold find_field.
  unfold proc_loc. 
  unfold e. Set Printing Depth 50. simpl. unfold load_value_of_type; simpl.
  (* b1 not change between m3 m8 *)
  generalize H6;intro.
  apply (Mem.load_alloc_other m3 0 (sizeof (Tpointer typ_SLv6_Processor))
    m8 b8 H25) in H6. 
  (* b1 not changed between m8 m10 *)
  (*apply load_store*)
Admitted.
*)

Lemma hasSPSR_true :
  forall m0 m0' m0'' e m vargs t m' v l b s em,
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m0'' ->
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    proc_state_related (of_mem proc m') e (Ok tt (mk_semstate l b s)) ->
    bool_val v T4 = Some true->
    Arm6_State.mode s = exn  em.
Proof.
Admitted.



Lemma hasSPSR_false :
  forall e m t m' v s,
    eval_expression (Genv.globalenv prog_adc) e m hasSPSR t m' v ->
    bool_val v T4 = Some false ->
    Arm6_State.mode s = usr.
Proof.
Admitted.

(*Lemma on proc_state_relates holds after copy_StatusRegister*)
Definition get_spsr :=
  Ecall (Evalof (Evar spsr T15) T15)
  (Econs (Evalof (Evar proc T3) T3)
    Enil) T8.

Axiom get_spsr_ok:
  forall e m t m' r,
    eval_expr (Genv.globalenv prog_adc) e m RV get_spsr t m' r ->
    m = m'.

Definition cp_SR :=
  Ecall
  (Evalof (Evar copy_StatusRegister T14) T14)
  (Econs
    (Eaddrof
      (Efield
        (Ederef (Evalof (Evar proc T3) T3) T6)
        cpsr T7) T8)
    (Econs
      (Ecall (Evalof (Evar spsr T15) T15)
        (Econs (Evalof (Evar proc T3) T3)
          Enil) T8) Enil)) T12.

Lemma same_cp_SR :
  forall e m l b s t m' v em,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    eval_expression (Genv.globalenv prog_adc) e m cp_SR t m' v ->
    (forall l b, proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b
      (Arm6_State.set_cpsr s (Arm6_State.spsr s em))))).
Proof.
  intros until em. intros psrel cpsr l' b'.
  inv cpsr. inv H. inv H4. inv H9. simpl in *.
  inv H5. inv H4. inv H5. inv H15. inv H4. inv H5.
  inv H14. inv H4. inv H3. inv H15. inv H5. inv H4. inv H5. inv H21.
  inv H13. simpl in *.
  (* Function spsr, get spsr from the current state *)
  apply (functions_behavior_ok e l b s vf0 fd0 m4 vargs0 t5 m2 vres0 l b s) 
    in psrel; [idtac|exact H18|exact H23].
  (* Function copy_StatusRegister, copy the current spsr to cpsr*)
  apply (functions_behavior_ok e l b s vf fd m2 vargs t3 m' vres l' b'
    (Arm6_State.set_cpsr s (Arm6_State.spsr s em)))
    in psrel; [idtac|exact H11|exact H16].
  exact psrel.
Qed.

(* Lemma on proc_state_relates holds after unpredictable*)
(* In fact, unpredictable in simlight is a annotation, which will print
   a error message. 
   For the moment, we consider it as a function call with an 
   empty body *)
Definition unpred :=
  Ecall
  (Evalof
    (Evar adc_compcert.unpredictable T16)
    T16) Enil T12.

Lemma same_unpred :
  forall e m s t m' v,
    proc_state_related (of_mem proc m) e (Ok tt s) ->
    eval_expression (Genv.globalenv prog_adc) e m unpred t m' v ->
    proc_state_related (of_mem proc m') e (Ko Arm6_Message.EmptyMessage).
Proof.
  intros until v. intros psrel unp.
  inv unp. inv H. inv H4. inv H9. inv H5.
  apply (funct_unpredictable e s vf fd m2 vargs t3 m' vres) in psrel;
  unfold unpredictable in psrel; unfold raise in psrel; 
  [exact psrel|exact H11|exact H16].
Qed.

(* Lemma on proc_state_relates holds after NZCV flag setting*)
Definition nflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef (Evalof (Evar proc T3) T3) T6)
      cpsr T7) N_flag T10)
  (Ecall (Evalof (Evar get_bit T17) T17)
    (Econs
      (Ecall (Evalof (Evar reg T2) T2)
        (Econs (Evalof (Evar proc T3) T3)
          (Econs 
            (Evalof (Evar d T4) T4) Enil))
        T1)
      (Econs (Eval (Vint (repr 31)) T9)
        Enil)) T10) T10.

Lemma same_nflag_assgnt :
  forall e m l b s d t m' v,
  proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
  d_func_related m e d ->
  eval_expression (Genv.globalenv prog_adc) e m nflag_assgnt t m' v->
  forall l b,
  proc_state_related (of_mem proc m') e
    (Ok tt
        (mk_semstate l b
           (Arm6_State.set_cpsr_bit s Nbit
              (Arm6_State.reg_content s d) [n31] )
         )
    ).
Proof.
Admitted.

Definition zflag_assgnt :=
  Eassign
  (Efield
    (Efield
      (Ederef 
        (Evalof (Evar proc T3) T3) T6)
      cpsr T7) Z_flag T10)
  (Econdition
    (Ebinop Oeq
      (Ecall (Evalof (Evar reg T2) T2)
        (Econs
          (Evalof (Evar proc T3) T3)
          (Econs
            (Evalof (Evar d T4) T4)
            Enil)) T1)
      (Eval (Vint (repr 0)) T9) T9)
    (Eval (Vint (repr 1)) T9)
    (Eval (Vint (repr 0)) T9) T9) T10.

Lemma same_zflag_assgnt :
  forall e m l b s d t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    d_func_related m e d ->
    eval_expression (Genv.globalenv prog_adc) e m zflag_assgnt t m' v->
    forall l b, proc_state_related (of_mem proc m') e 
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Zbit
        (if Util.zeq (Arm6_State.reg_content s d) 0
         then repr 1
         else repr 0)))).
Proof.
Admitted.

Definition cflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef
        (Evalof (Evar proc T3) T3)
        T6) cpsr T7) C_flag T10)
  (Ecall
    (Evalof 
      (Evar CarryFrom_add3 T18) T18)
    (Econs
      (Evalof (Evar old_Rn T1) T1)
      (Econs
        (Evalof
          (Evar shifter_operand T1)
          T1)
        (Econs
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T10)
            T10) Enil))) T10) T10.

Lemma same_cflag_assgnt:
  forall m e l b s0 s n so t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    n_func_related m e n ->
    so_func_related m e so ->
    eval_expression (Genv.globalenv prog_adc) e m cflag_assgnt t m' v->
    forall l b, proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Cbit
        (Arm6_Functions.CarryFrom_add3 (Arm6_State.reg_content s0 n) so
          (Arm6_State.cpsr (st (mk_semstate l b s))) [Cbit])))).
Proof.
Admitted.

Definition vflag_assgnt:=
  Eassign
  (Efield
    (Efield
      (Ederef
        (Evalof (Evar proc T3) T3)
        T6) cpsr T7) V_flag T10)
  (Ecall
    (Evalof
      (Evar OverflowFrom_add3 T19)
      T19)
    (Econs
      (Evalof (Evar old_Rn T1) T1)
      (Econs
        (Evalof
          (Evar shifter_operand T1)
          T1)
        (Econs
          (Evalof
            (Efield
              (Efield
                (Ederef
                  (Evalof (Evar proc T3) T3)
                  T6) cpsr T7) C_flag T10)
            T10) Enil))) T10) T10.

Lemma same_vflag_assgnt:
  forall m e l b s0 s n so t m' v,
    proc_state_related (of_mem proc m) e (Ok tt (mk_semstate l b s)) ->
    n_func_related m e n ->
    so_func_related m e so ->
    eval_expression (Genv.globalenv prog_adc) e m vflag_assgnt t m' v->
    proc_state_related (of_mem proc m') e
      (Ok tt (mk_semstate l b (Arm6_State.set_cpsr_bit s Arm6_SCC.Vbit
        (Arm6_Functions.OverflowFrom_add3 (Arm6_State.reg_content s0 n) so
           (Arm6_State.cpsr (st (mk_semstate l b s))) [Cbit])))).
Proof.
Admitted.


(* During function execution, none other parameters are changed*)
Lemma cp_SR_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m cp_SR Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma reg_S_not_changed :
  forall e m vargs t m' v,
    eval_funcall (Genv.globalenv prog_adc) m (Internal fun_internal_reg) 
    vargs t m' v ->
    param_val S m e = param_val S m' e.
Proof.
Admitted.

Lemma reg_mem_not_changed:
  forall m vargs t m' v,
    eval_funcall (Genv.globalenv prog_adc) m (Internal fun_internal_reg) 
    vargs t m' v ->
    m = m'.
Proof.
  intros until v. intro ef.
  inv ef.
Admitted. 


Lemma rn_ass_S_not_changed:
  forall m0 m0' vargs m e v m', 
    alloc_variables empty_env m0 
      (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m0' ->
    bind_parameters e m0' fun_internal_ADC.(fn_params) vargs m ->
    list_norepet 
    (var_names fun_internal_ADC.(fn_params) ++ var_names fun_internal_ADC.(fn_vars)) ->
    eval_expression (Genv.globalenv prog_adc) e m oldrn_assgnt Events.E0 m' v ->
    param_val S m e = param_val S m' e.
Proof.
  intros until m'. intros av bp ln evex.
  inv_alloc_vars e.
  pose(e:=
    (PTree.set old_Rn (b6, Tint I32 Unsigned)
      (PTree.set shifter_operand (b5, Tint I32 Unsigned)
        (PTree.set n (b4, Tint I8 Unsigned)
          (PTree.set d (b3, Tint I8 Unsigned)
            (PTree.set cond (b2, Tint I32 Signed)
              (PTree.set S (b0, Tint I8 Signed)
                (PTree.set proc (b1, Tpointer typ_SLv6_Processor)
                  empty_env))))))));
  fold e in bp, evex |-*.
  inv_bind_params m.
  repeat rrw_block.
  unfold store_value_of_type in *;simpl in str,str0,str1,str2,str3,str4.
  
  (* begin with assgn expr *)
  (* eval_expression from m to m'*)
  inv evex. 
  (* eval assignment, left:m->m13, right:m13->14, storage of Rn:m14->m' *)
  inv H. 
  (* esr_rval in m' *)
  inv H0.
  simpl in H11.
  (* eval Evar from m to m13, m=m13 *)
  inv H5. 
  (* eval Ecall from m13 to m14 *)  
  inv H6. 
  (* eval Evalof from m13 to m1 *)
  inv H2.
  (* eval Evar, m13=m1*)
  inv H13.
  (* first param of reg, proc *)
  (* eval_exprlist from m1 to m15 *)
  inv H3.
  (* eval Evalof from m1 to m13*)
  inv H6.
  (* eval Evar m1=m13*)
  inv H3.
  (* second param of reg, n *)
  (* eval_exprlist from m13 to m15 *)
  inv H19.
  (* eval Evalof from m13 to m1 *)
  inv H3.
  (* eval Evar m13=m1*)
  inv H6.
  (* no more param *)
  inv H18.
  (* function fd is reg *)
  injection H9;intros Hres Hargs;subst;clear H9 H17.
  inv H5.
  (* esl_var_global in m15 *)
  inv H1;[discriminate|].
  unfold Genv.find_symbol in H5;simpl in H5.
  (* b7=-5*)
  injection H5;intro;subst;clear H2 H5 H14.
  (* vf = Vptr (-5) w0 *)
  unfold load_value_of_type in H6;simpl in H6;injection H6;intro;subst;clear H6.
  rewrite Genv.find_funct_find_funct_ptr in H16.
  injection H16;intro Hfd;rewrite<-Hfd in *;clear Hfd fd H16.
  (* eval_funcall reg from m15 to m14*)
  inv H21.
  (* exec_stmt from m13 to m16 *)
  inv H5. simpl in H6.
  (* eval_expression reg_m from m13 to m16 *)
  inv H16.
  (* eval Ecall reg_m from m13 to m16 *)
  inv H.
  (* eval Evalof from m13 to m17 *)
  inv H17.
  (* eval Evar m13 = m17 *)
  inv H22.
  (* eval_exprlist from m17 to m18 *)
  inv H18.
  (* first param of reg_m, proc *)
  (* eval Evalof from m17 to m13 *)
  inv H17.
  (* eval Evar m17=m13 *)
  inv H18.
  (* second param of reg_m, reg_id *)
  inv H27.
  (* eval evalof from m13 to m17 *)
  inv H17.
  (* eval evar m13=m17*)
  inv H18.
  (* third param of reg_m, proc->cpsr *)
  inv H26.
  (* eval Evalof from m17 to m13*)
  inv H17.
  (* eval Efield from m17 yo m13*)
  inv H18.
  (* eval Efield from m17 to m13*)
  inv H28.
  (* eval Ederef from m17 to m13*)
  inv H26.
  (* eval Evalof from m17 to m13*)
  inv H17.
  (* eval Evar m17=m13*)
  inv H18.
  (* no more param for reg_m,m13=m18*)
  inv H27.
  (* v7 = Eval vres0 T1*)
  inv H5.
  (* esr_valof in m18, find reg_m in golbal *)
  inv H19.
  (* e0 *)
  inv_alloc_vars e0.
  pose(e0:=(PTree.set adc_compcert.reg_id (b9, Tint I8 Unsigned)
    (PTree.set proc (b8, Tpointer typ_SLv6_Processor) empty_env)));
  fold e0 in H13,H20,H2,H9.
  (* esl_var_global in m18 *)
  inv H9;[discriminate|].
  (* find the value of b7 *)
  injection H16;intro;rewrite<-H in *;clear H H16 b7.
  unfold load_value_of_type in H17;simpl in H17.
  injection H17;intro;rewrite<-H in *;clear H17 H22 H vf.
  rewrite Genv.find_funct_find_funct_ptr in H24.
  injection H24;intro;rewrite<-H in *;clear H H24 fd.
  (* eval_funcall reg_m from m18 to m16*)
  inv H29.
  (* exec_stmt of reg_m from m19 to m20 *)
  inv H17.
  simpl in H18.
  (* eval_expression from m19 to m20*)
  inv H24.
  (* eval evalof from m19 to m20*)
  inv H.
  (* eval Ederef from m19 to m20*)
  inv H27.
  (* *)
Admitted.





  

(*
  (* reg is in loc env *)
  assert (reg_not_loc: e!reg = None).
  unfold e. simpl. reflexivity.
  inv H5. inv H1. rewrite reg_not_loc in H9. discriminate H9. clear H3.

  (* ofs is w0 *)
  inv H5. clear H2. inv H6. inv H16.
  destruct eq_dec; [idtac|discriminate H0]. clear e0. inv H0.

  (*
  (* open internal function reg *)
  inv H21. inv H1. inv H20. inv H21.
*)


  (* nextblock is not change from Mem.store on memory *)
  generalize alc12; intro.
  apply Mem.valid_new_block in alc1. unfold Mem.valid_block in alc1.
  apply Mem.nextblock_store in st0.
  apply Mem.nextblock_store in st2.
  apply Mem.nextblock_store in st3.
  apply Mem.nextblock_store in st4.
  apply Mem.nextblock_store in st5.
  apply Mem.nextblock_store in st6.
  rewrite <- st6 in st5. rewrite <- st5 in st4. rewrite <- st4 in st3. 
  rewrite <- st3 in st2. rewrite <- st2 in st0.
  rewrite <- st0 in alc1.

  (* b0 < b6 *)
  generalize H19; intros.
  apply Mem.alloc_result in H19. rewrite <- H19 in alc1.
  apply (Zlt_trans b4) in alc1; [idtac|exact lt411]. 
  apply (Zlt_trans b0) in alc1; [idtac|exact lt0].

  (* expand bind_parameters *)
  inv H2. inv H23. inv H24. simpl in H16, H15.
  inversion H16. rewrite <- H2 in *. clear b8 H16 H2.
  inversion H15. rewrite H2 in *. clear b7 H15 H2.

  (* between m15 and m17 *)  
  assert (load_value_of_type (Tint I8 Unsigned) m17 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m15 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_alloc_unchanged m15 0 
    (sizeof (Tpointer typ_SLv6_Processor)) m17 (Mem.nextblock m15));
  [exact H1|unfold Mem.valid_block; exact alc1].
  
  (* between m17 and m1 *)
  generalize H18; intro.
  apply Mem.valid_new_block in H1. unfold Mem.valid_block in H1.
  apply Mem.alloc_result in H18.
  apply (Zlt_trans b0) in H1; [idtac|exact alc1].
  assert (load_value_of_type (Tint I8 Unsigned) m1 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m17 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_alloc_unchanged m17 0 
    (sizeof (Tint I8 Unsigned)) m1 b6);
  [exact H2|unfold Mem.valid_block; exact H1].
  rewrite <- H6 in H. clear H6.

  (* between m1 and m18 *)
  unfold store_value_of_type in H22, H21; simpl in H22, H21.
  assert (load_value_of_type (Tint I8 Unsigned) m18 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m1 b0 w0). 
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m1 ((Mem.nextblock m15)) (signed w0) v7);
    [exact H22|left;apply Zlt_not_eq in alc1; exact alc1].
  rewrite <- H6 in H. clear H6.

  (* betwwen m18 and m13 *)
  assert (load_value_of_type (Tint I8 Unsigned) m13 b0 w0 =
  load_value_of_type (Tint I8 Unsigned) m18 b0 w0). 
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint8unsigned m18 b6 (signed w0) v8);
    [exact H21|left; apply Zlt_not_eq in H1; rewrite <- H18 in H1; exact H1].
  rewrite <- H6 in H. clear H6.

  (* between m13 and m16 *)
  pose (e0 := (PTree.set adc_compcert.reg_id (b6, Tint I8 Unsigned)
            (PTree.set proc (Mem.nextblock m15, Tpointer typ_SLv6_Processor)
               empty_env))).
  (*fold e0 in H3.
  inv H3. inv H15.*)
  inv H3. fold e0 in H15. inv H15.  inv H3. inv H16.


  apply (reg_S_not_changed e m15 vargs t3 m14 v6) in H21.
  unfold param_val in H21. unfold e in H21; simpl in H21.
  unfold store_value_of_type in H12; simpl in H12.

  assert (Heqm'm14: load_value_of_type (Tint I8 Signed) m' b0 w0=
  load_value_of_type (Tint I8 Signed) m14 b0 w0).
  unfold load_value_of_type; simpl.
  apply (Mem.load_store_other AST.Mint32 m14 b5 (unsigned ofs) v). exact H12.
  left.
  inv H7; [idtac|inv H2]. 
  unfold e in H3; simpl in H3. inversion H3. rewrite <- H0 in *.
  clear b5 H0.
  apply (diff_block m11 (sizeof (Tint I32 Unsigned)) b4) in alc12;
    [apply (Zlt_trans b0) in alc12; 
      [apply Zlt_not_eq in alc12; exact alc12|exact lt0] |exact alc11].
  
  rewrite H21. rewrite Heqm'm14. reflexivity.
Qed.
*)

Lemma rn_ass_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m oldrn_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma set_reg_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m set_regpc Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma unpred_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m unpred Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma nf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m nflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma zf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m zflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma vf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m vflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma cf_params_not_changed:
  forall m e v m' i, 
    eval_expression (Genv.globalenv prog_adc) e m cflag_assgnt Events.E0 m' v ->
    param_val i m e = param_val i m' e.
Proof.
Admitted.

Lemma same_bool : forall b, b&&b = b.
Proof.
  destruct b;simpl;reflexivity.
Qed.

Theorem related_aft_ADC: forall e m0 m1 m2 mfin vargs s out sbit cond d n so,
  alloc_variables empty_env m0 (fun_internal_ADC.(fn_params) ++ fun_internal_ADC.(fn_vars)) e m1 ->
  bind_parameters e m1 fun_internal_ADC.(fn_params) vargs m2 ->
(* TODO: valid_access needs to be more precise *)
  (forall m ch b ofs, Mem.valid_access m ch b ofs Readable) ->
  proc_state_related (of_mem proc m2) e (Ok tt (mk_semstate nil true s)) ->
  sbit_func_related m2 e sbit ->
  cond_func_related m2 e cond ->
  d_func_related m2 e d ->
  n_func_related m2 e n ->
  so_func_related m2 e so ->
(* Comparison between eval_funcall, exec_stmt:
   [eval_funcall] is big step semantic. It can be seen as 6 steps, 
   and we can observe 4 times of memory changes.
   1. Check there are no repetitive parameters in function parameter list;
   2. Allocate function parameters into memory and fill them in the empty local environment (m0->m1);
   3. Bind these parameters with there initial values (m1->m2);
   4. Execute all the statement of the function body (m2->m3);
   5. Clean up the memory which are used to store the local parameters when
   execution finishes (m3->m4).
   This final memory doesn't contain the final [proc] we expect. It is in [m3], but in [m4],
   their memory blocks are freed.
   [exec_stmt] is also big step semantic. It indicates the outcome of 
   statement execution [Out_break], [Out_continue], [Out_normal] and [Out_return].
   The final memory state is the memory which contains the final values of parameters.
   The final [proc] is in this memory state which we want to relate.*)
  exec_stmt (Genv.globalenv prog_adc) e m2 fun_internal_ADC.(fn_body) Events.E0 mfin out ->
  proc_state_related (of_mem proc mfin) e (S.ADC_step sbit cond d n so (mk_semstate nil true s)). 
Proof.
  
  intros until so.
  intros al bi valacc psrel sfrel cfrel dfrel nfrel sofrel exstmt.

  (* expand the whole statement of ADC, from m2 to mfin *)
  inv exstmt; [idtac | nod];
  apply Events.Eapp_E0_inv in H3; destruct H3; subst.
  rename H4 into rn_assgnt, H7 into main_p.
  (* Old_Rn assignment, from m2 to m3 *)
  inv rn_assgnt;
  rename H2 into rn_assgnt.
  (* the projection relation between state and other parameters
     still hold after execute old_rn assignment, from m2 to m3 *)
  apply (oldrn_assgnt_ok e m2 nil true s Events.E0 m3 v) in psrel; 
    [idtac|exact rn_assgnt].
  unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 S) in sfrel;
    [idtac | exact rn_assgnt];
  fold (bit_proj m3 e S) in sfrel; fold (sbit_func_related m3 e sbit) in sfrel.
  unfold cond_func_related in cfrel; unfold cond_proj in cfrel.
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert.cond) in cfrel;
    [idtac | exact rn_assgnt];
  fold (cond_proj m3 e) in cfrel; fold (cond_func_related m3 e cond) in cfrel.
  unfold d_func_related in dfrel; unfold reg_proj in dfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert.d) in dfrel;
    [idtac | exact rn_assgnt];
  fold (reg_proj m3 e adc_compcert.d) in dfrel; fold (d_func_related m3 e d) in dfrel.
  unfold n_func_related in nfrel; unfold reg_proj in nfrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 adc_compcert.n) in nfrel;
    [idtac | exact rn_assgnt]; 
  fold (reg_proj m3 e adc_compcert.n) in nfrel; fold (n_func_related m3 e n) in nfrel.
  unfold so_func_related in sofrel; unfold bits_proj in sofrel;
  rewrite (rn_ass_params_not_changed m2 e v m3 shifter_operand) in sofrel;
    [clear rn_assgnt | exact rn_assgnt];
  fold (bits_proj m3 e shifter_operand) in sofrel;
  fold (so_func_related m3 e so) in sofrel.
  (* ConditionPassed, from m3 to m4, m3 = m4 *)
  inv main_p;
  rename H5 into condpass, H8 into cp_b, H9 into main_p, H4 into evs;
  generalize condpass;intro condpass';
      simpl in cp_b;
      apply Events.Eapp_E0_inv in evs; destruct evs; subst;
      apply no_effect_condpass in condpass0;
      rewrite condpass0 in *;clear condpass0.
      (* ConditionPassed(&proc->cpsr, cond) has the same value as 
         Arm6_Functions.State.ConditionPassed s cond, in m4 *)
      apply (condpass_bool m0 m1 e m4 Events.E0 m4 v1 cond s) in cp_b;
        [idtac| exact al| exact condpass'].
      (* two cases, the boolean value of ConditionPassed *)
      destruct b.
        (* ConditionPassed(&proc->cpsr, cond) evaluates to true *)
        (* set_reg_or_pc, from m4 to m5 *)
        inv main_p; [idtac | nod];
        rename H4 into setreg, H7 into main_p, H3 into evs;
        apply Events.Eapp_E0_inv in evs; destruct evs; subst.
        (* projection relation between state and other parameters after execute
           set_reg_or_pc, from m4 to m5 *)
        inv setreg;
        rename H2 into setreg;
        apply (same_setregpc e m4 nil true s s Events.E0 m5 v0 d n so) 
        with nil (Util.zne d 15) in psrel;
          [idtac | fold set_regpc in setreg; apply setreg].
        unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
        rewrite (set_reg_params_not_changed m4 e v0 m5 S) in sfrel;
          [idtac | exact setreg];
        fold (bit_proj m5 e S) in sfrel; fold (sbit_func_related m5 e sbit) in sfrel.
        unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
        rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert.cond) in cfrel;
          [idtac | exact setreg];
        fold (cond_proj m5 e) in cfrel; fold (cond_func_related m5 e cond) in cfrel.
        unfold d_func_related in dfrel; unfold reg_proj in dfrel;
        rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert.d) in dfrel;
          [idtac | exact setreg];
        fold (reg_proj m5 e adc_compcert.d) in dfrel; 
        fold (d_func_related m5 e d) in dfrel.
        unfold n_func_related in nfrel; unfold reg_proj in nfrel;
        rewrite (set_reg_params_not_changed m4 e v0 m5 adc_compcert.n) in nfrel;
          [idtac | exact setreg]; 
        fold (reg_proj m5 e adc_compcert.n) in nfrel;
        fold (n_func_related m5 e n) in nfrel.
        unfold so_func_related in sofrel; unfold bits_proj in sofrel;
        rewrite (set_reg_params_not_changed m4 e v0 m5 shifter_operand) in sofrel;
          [clear setreg | exact setreg];
        fold (bits_proj m5 e shifter_operand) in sofrel;
        fold (so_func_related m5 e so) in sofrel.
        (* S == 1 && d == 15, from m5 to m6, has no effect on memory, m5 = m6 *)
        inv main_p;
          rename H5 into sd, H8 into sd_b, H9 into main_p, H4 into evs;
          generalize sd;intro sd';
          simpl in sd_b;
          apply no_effect_is_S_set_and_is_pc in sd;
          rewrite sd in *;clear sd;
          apply Events.Eapp_E0_inv in evs; destruct evs; subst.
        (* S == 1 && d == 15 has the same value as in Coq side, in m6 *)
        apply (S_pc_bool e m6 Events.E0 m6 v2 sbit d) in sd_b;
        [idtac|exact sfrel|exact dfrel|exact sd'].
        (* two cases on the boolean value of S == 1 && d == 15 *)
        destruct b.
          (* ((S == 1) && (d == 15)) evaluates to true *)
          (* CurrentModeHasSPSR has no effect on memory, from m6 to m7, m6=m7 *)
          inv main_p;
          rename H5 into hasspsr, H8 into spsr_b, H9 into main_p, H4 into evs;
          generalize hasspsr;intro hasspsr1;
            simpl in spsr_b;
            apply Events.Eapp_E0_inv in evs; destruct evs; subst.
            apply if_hasSPSR_ok in hasspsr;
            rewrite hasspsr in *;clear hasspsr.
          (* two cases on the boolean value of CurrentModeHasSPSR *)
          destruct b.
            (* CurrentModeHasSPSR evaluate to true *)
            apply (hasSPSR_true m0 m1 m2 e m7 vargs Events.E0 m7 v3
              nil (Util.zne d 15)
              (Arm6_State.set_reg s d
                (add (add (Arm6_State.reg_content s n) so)
                  (Arm6_State.cpsr s) [Cbit])) und) in spsr_b;
            [idtac |exact al|exact bi|exact hasspsr1|exact psrel].
            (* copy_StatusRegister, from m7 to mfin *)
            inv main_p;
            rename H2 into cp_sr.
            (*generalize psrel; intro psrelm7.*)
            (* projection relation between state and other parameters still hold
               after executing copy_StatusRegister, from m7 to mfin.
               And finally get the projection relation on memory mfin *)
            apply (same_cp_SR e m7 nil (Util.zne d 15) 
              (Arm6_State.set_reg s d
                (add (add (Arm6_State.reg_content s n) so)
                  (Arm6_State.cpsr s) [Cbit])) Events.E0 mfin v4 und) 
            with nil (Util.zne d 15) in psrel;
              [idtac | exact cp_sr ].
            unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
            rewrite (cp_SR_params_not_changed m7 e v4 mfin S) in sfrel;
              [idtac | exact cp_sr];
            fold (bit_proj mfin e S) in sfrel;
            fold (sbit_func_related mfin e sbit) in sfrel.
            unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
            rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert.cond) 
              in cfrel;
              [idtac | exact cp_sr];
            fold (cond_proj mfin e) in cfrel;
            fold (cond_func_related mfin e cond) in cfrel.
            unfold d_func_related in dfrel; unfold reg_proj in dfrel;
            rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert.d) in dfrel;
              [idtac | exact cp_sr];
            fold (reg_proj mfin e adc_compcert.d) in dfrel;
            fold (d_func_related mfin e d) in dfrel.
            unfold n_func_related in nfrel; unfold reg_proj in nfrel;
            rewrite (cp_SR_params_not_changed m7 e v4 mfin adc_compcert.n) in nfrel;
              [idtac | exact cp_sr]; 
            fold (reg_proj mfin e adc_compcert.n) in nfrel;
            fold (n_func_related mfin e n) in nfrel.
            unfold so_func_related in sofrel; unfold bits_proj in sofrel;
            rewrite (cp_SR_params_not_changed m7 e v4 mfin shifter_operand) in sofrel;
              [clear cp_sr | exact cp_sr];
            fold (bits_proj mfin e shifter_operand) in sofrel;
            fold (so_func_related mfin e so) in sofrel.
            (* expand ADC_step *)
            unfold S.ADC_step; unfold _get_st; unfold bind_s;
            unfold bind; simpl.
            rewrite cp_b;rewrite sd_b; simpl.
            unfold if_CurrentModeHasSPSR; unfold block; unfold fold_left;
            unfold _get_bo; unfold bind_s; unfold next; unfold bind; simpl;
            unfold _Arm_State.set_reg.
            rewrite spsr_b; simpl; unfold _Arm_State.set_reg. 
            unfold _Arm_State.set_cpsr;
            unfold _set_bo; unfold ok_semstate; unfold loc; unfold st. 
            rewrite same_bool.
            (* The same projection relation as the one in hypothesis *)
            exact psrel.
            
            (* CurrentModeHasSPSR(proc) evaluates to false *)
            apply (hasSPSR_false e m7 Events.E0 m7 v3
              (Arm6_State.set_reg s d
                (add (add (Arm6_State.reg_content s n) so)
                  (Arm6_State.cpsr s) [Cbit]))) in spsr_b;
            [idtac |exact hasspsr1].
            (* meet unpredictable *)
            inv main_p; rename H2 into unp.
            (* projection relation between state and other parameters still hold
               after unpredictable, from m7 to mfin.*)
            apply (same_unpred e m7 
              (mk_semstate nil (Util.zne d 15) (Arm6_State.set_reg s d
                (add (add (Arm6_State.reg_content s n) so)
                  (Arm6_State.cpsr s) [Cbit]))) Events.E0 mfin v4) in psrel;
            [idtac | exact unp].
            unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
            rewrite (unpred_params_not_changed m7 e v4 mfin S) in sfrel;
              [idtac | exact unp];
            fold (bit_proj mfin e S) in sfrel; 
            fold (sbit_func_related mfin e sbit) in sfrel.
            unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
            rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert.cond) 
              in cfrel;
              [idtac | exact unp];
            fold (cond_proj mfin e) in cfrel;
            fold (cond_func_related mfin e cond) in cfrel.
            unfold d_func_related in dfrel; unfold reg_proj in dfrel;
            rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert.d) 
              in dfrel;
              [idtac | exact unp];
            fold (reg_proj mfin e adc_compcert.d) in dfrel;
            fold (d_func_related mfin e d) in dfrel.
            unfold n_func_related in nfrel; unfold reg_proj in nfrel;
            rewrite (unpred_params_not_changed m7 e v4 mfin adc_compcert.n) in nfrel;
              [idtac | exact unp]; 
            fold (reg_proj mfin e adc_compcert.n) in nfrel;
            fold (n_func_related mfin e n) in nfrel.
            unfold so_func_related in sofrel; unfold bits_proj in sofrel;
            rewrite (unpred_params_not_changed m7 e v4 mfin shifter_operand) 
              in sofrel;
              [clear unp | exact unp];
            fold (bits_proj mfin e shifter_operand) in sofrel;
            fold (so_func_related mfin e so) in sofrel.
            (* expand ADC_step *)
            unfold S.ADC_step; unfold _get_st; unfold bind_s;
            unfold bind; simpl.
            rewrite cp_b; rewrite sd_b; simpl.
            unfold if_CurrentModeHasSPSR; unfold block; unfold fold_left;
            unfold _get_bo; unfold bind_s; unfold next; unfold bind;
            simpl; unfold _Arm_State.set_reg.
            rewrite spsr_b; simpl.
            (* The same projection relation as the one in hypothesis *)
            exact psrel.
          (* ((S == 1) && (d == 15)) evaluates to false *)
          (* S==1 has no effect on memory m6 = m7 *)
          inv main_p;
          rename H5 into is_s, H8 into s_b, H9 into main_p, H4 into evs;
          generalize is_s;intros is_s';
            simpl in s_b; 
            apply no_effect_is_S_set in is_s;
            rewrite is_s in *;clear is_s;
            apply Events.Eapp_E0_inv in evs; destruct evs; subst.
          (* S==1 has the same result as in Coq in m7 *)
          apply (S_bool m0 e m1 m7 Events.E0 m7 v3 sbit) in s_b;
            [idtac|exact al|exact sfrel|exact is_s'].
          (* two cases on the bool value of S==1 *)
          destruct b.
            (* S == 1 evaluates to true *)
            (* N_flag assignment from m7 to m8 *)
            inv main_p ;[idtac | nod];
            rename H4 into nf, H7 into main_p, H3 into evs;
            apply Events.Eapp_E0_inv in evs; destruct evs; subst.
            (* projection relation between state and other parameters still hold
               after N_flag assignment, from m7 to m8 *)
            inv nf; rename H2 into nf;
            pose (s0 :=  Arm6_State.set_reg s d
                       (add (add (Arm6_State.reg_content s n) so)
                          (Arm6_State.cpsr s) [Cbit]));
            fold s0 in psrel.
            eapply (same_nflag_assgnt e m7 nil (Util.zne d 15)
              s0 d Events.E0 m8 v4) in psrel;
            [idtac | exact dfrel | exact nf].
            unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
            rewrite (nf_params_not_changed m7 e v4 m8 S) in sfrel;
              [idtac | exact nf];
            fold (bit_proj m8 e S) in sfrel;
            fold (sbit_func_related m8 e sbit) in sfrel.
            unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
            rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert.cond) in cfrel;
              [idtac | exact nf];
            fold (cond_proj m8 e) in cfrel;
            fold (cond_func_related m8 e cond) in cfrel.
            unfold d_func_related in dfrel; unfold reg_proj in dfrel;
            rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert.d) in dfrel;
              [idtac | exact nf];
            fold (reg_proj m8 e adc_compcert.d) in dfrel;
            fold (d_func_related m8 e d) in dfrel.
            unfold n_func_related in nfrel; unfold reg_proj in nfrel;
            rewrite (nf_params_not_changed m7 e v4 m8 adc_compcert.n) in nfrel;
              [idtac | exact nf]; 
            fold (reg_proj m8 e adc_compcert.n) in nfrel;
            fold (n_func_related m8 e n) in nfrel.
            unfold so_func_related in sofrel; unfold bits_proj in sofrel;
            rewrite (nf_params_not_changed m7 e v4 m8 shifter_operand) in sofrel;
              [clear nf | exact nf];
            fold (bits_proj m8 e shifter_operand) in sofrel;
            fold (so_func_related m8 e so) in sofrel.
            (* Z_flag assignment from m8 to m9 *)
            inv main_p ;[idtac | nod];
            rename H4 into zf, H7 into main_p, H3 into evs;
            apply Events.Eapp_E0_inv in evs; destruct evs; subst.
            (* projection relation between state and other parameters still hold
               after Z_flag assignment, from m8 to m9 *)
            inv zf; rename H2 into zf;
            pose (s1 := Arm6_State.set_cpsr_bit s0 Nbit
              (Arm6_State.reg_content s0 d) [n31]);
            revert psrel; fold s1; intro psrel;
            eapply (same_zflag_assgnt e m8 nil (Util.zne d 15) s1
              d Events.E0 m9 v5) in psrel;
            [idtac| exact dfrel | exact zf].
            unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
            rewrite (zf_params_not_changed m8 e v5 m9 S) in sfrel;
              [idtac | exact zf];
            fold (bit_proj m9 e S) in sfrel;
            fold (sbit_func_related m9 e sbit) in sfrel.
            unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
            rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert.cond) in cfrel;
              [idtac | exact zf];
            fold (cond_proj m9 e) in cfrel;
            fold (cond_func_related m9 e cond) in cfrel.
            unfold d_func_related in dfrel; unfold reg_proj in dfrel;
            rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert.d) in dfrel;
              [idtac | exact zf];
            fold (reg_proj m9 e adc_compcert.d) in dfrel;
            fold (d_func_related m9 e d) in dfrel.
            unfold n_func_related in nfrel; unfold reg_proj in nfrel;
            rewrite (zf_params_not_changed m8 e v5 m9 adc_compcert.n) in nfrel;
              [idtac | exact zf]; 
            fold (reg_proj m9 e adc_compcert.n) in nfrel;
            fold (n_func_related m9 e n) in nfrel.
            unfold so_func_related in sofrel; unfold bits_proj in sofrel;
            rewrite (zf_params_not_changed m8 e v5 m9 shifter_operand) in sofrel;
              [clear zf | exact zf];
            fold (bits_proj m9 e shifter_operand) in sofrel; 
            fold (so_func_related m9 e so) in sofrel.
            (* C_flag assignment from m9 to m10 *)
            inv main_p ;[idtac | nod];
            rename H4 into cf, H7 into vf, H3 into evs;
            apply Events.Eapp_E0_inv in evs; destruct evs; subst.
            (* projection relation between state and other parameters still hold
               after C_flag assignment, from m9 to m10 *)
            inv cf; rename H2 into cf;
            pose (s2 := Arm6_State.set_cpsr_bit s1 Zbit
              (if Util.zeq (Arm6_State.reg_content s1 d) 0
                then repr 1
                else repr 0));
            revert psrel; fold s2; intro psrel;
            eapply (same_cflag_assgnt m9 e nil (Util.zne d 15) s s2
              n so Events.E0 m10 v6) in psrel;
            [idtac| exact nfrel | exact sofrel| exact cf]. 
            unfold sbit_func_related in sfrel; unfold bit_proj in sfrel;   
            rewrite (cf_params_not_changed m9 e v6 m10 S) in sfrel;
              [idtac | exact cf];
            fold (bit_proj m10 e S) in sfrel;
            fold (sbit_func_related m10 e sbit) in sfrel.
            unfold cond_func_related in cfrel; unfold cond_proj in cfrel;
            rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert.cond) in cfrel;
              [idtac | exact cf];
            fold (cond_proj m10 e) in cfrel;
            fold (cond_func_related m10 e cond) in cfrel.
            unfold d_func_related in dfrel; unfold reg_proj in dfrel;
            rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert.d) in dfrel;
              [idtac | exact cf];
            fold (reg_proj m10 e adc_compcert.d) in dfrel;
            fold (d_func_related m10 e d) in dfrel.
            unfold n_func_related in nfrel; unfold reg_proj in nfrel;
            rewrite (cf_params_not_changed m9 e v6 m10 adc_compcert.n) in nfrel;
              [idtac | exact cf]; 
            fold (reg_proj m10 e adc_compcert.n) in nfrel;
            fold (n_func_related m10 e n) in nfrel.
            unfold so_func_related in sofrel; unfold bits_proj in sofrel;
            rewrite (cf_params_not_changed m9 e v6 m10 shifter_operand) in sofrel;
              [clear cf | exact cf];
            fold (bits_proj m10 e shifter_operand) in sofrel;
            fold (so_func_related m10 e so) in sofrel.
            (* projection relation between state still hold
               after V_flag assignment, from m10 to mfin *)
            unfold st in psrel.
            inv vf; rename H2 into vf;
            pose (s3 := Arm6_State.set_cpsr_bit s2 Cbit
              (Arm6_Functions.CarryFrom_add3
                (Arm6_State.reg_content s n) so
                (Arm6_State.cpsr s2) [Cbit]));
            revert psrel; fold s3; intro psrel;
            eapply (same_vflag_assgnt m10 e nil (Util.zne d 15) s s3
              n so Events.E0 mfin v7) in psrel;
            [clear vf| exact nfrel | exact sofrel| exact vf].
            (* expand ADC_step, simplifiy all the if else case *)
            unfold S.ADC_step; unfold _get_st; unfold bind_s; unfold bind; simpl.
            rewrite cp_b; simpl. 
            unfold block; unfold fold_left at 1; unfold next; 
            unfold bind at 1 2; unfold _get_bo at 1;
            unfold bind_s at 1; unfold bind at 1; unfold bind at 1; 
            unfold set_reg; simpl; unfold _Arm_State.set_reg. 
            fold s0.
            rewrite sd_b; rewrite s_b; simpl.
            (* Nflag *)
            unfold bind at 5. unfold _get_bo at 2. unfold bind_s at 1. 
            unfold bind at 5. unfold bind at 5.
            simpl; unfold _Arm_State.set_cpsr_bit at 1. 
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            unfold _set_bo at 1.  simpl. unfold ok_semstate.
            (* Zflag *)
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
            (* Cflag *)
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
            (* Vflag *)
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            unfold bind at 5. simpl; unfold _Arm_State.set_cpsr_bit at 1.
            unfold _get_bo at 2. unfold bind_s at 1. unfold bind at 5.
            simpl. unfold _set_bo at 1. simpl. unfold ok_semstate.
            unfold bind at 4. unfold loc at 1. unfold bo at 1. unfold bo at 3.
            unfold st at 1. unfold st at 3.
            unfold bind at 3. unfold loc at 1. unfold bo at 1. unfold bo at 5.
            unfold st at 1. unfold st at 5.
            unfold bind at 2. unfold loc at 1. unfold bo at 1. unfold bo at 9.
            unfold st at 1. unfold st at 9.
            (* simplify the bo and st of semstate *)
            unfold bind at 1. unfold _get_bo at 2. unfold bind_s at 1.
            unfold bind at 1. unfold bo at 1.
            unfold _set_bo at 1. unfold loc at 1. unfold st at 1.
            unfold ok_semstate.
            unfold _get_bo at 1. unfold bind_s at 1. unfold bind at 1.
            unfold loc at 1. unfold bo. unfold st at 1. unfold st.
            fold s1. fold s2. fold s3. unfold st in psrel.
            rewrite same_bool; rewrite same_bool; rewrite same_bool;
            rewrite same_bool; rewrite same_bool.
            (* get the same projection relation as the one in hypothesis *)
            exact psrel.
            (* S == 1 evaluates to false *)
            (* Skip statement from m7 to mfin, m7 = mfin *)
            inv main_p.
            (* expand ADC_step *)
            unfold S.ADC_step; unfold _get_st; unfold bind_s; unfold bind; simpl.
            rewrite cp_b; rewrite sd_b; rewrite s_b; simpl.
            unfold block. unfold fold_left. unfold next.
            unfold bind at 3. simpl; unfold _Arm_State.set_reg.
            unfold _get_bo at 2. unfold bind_s at 1. unfold _set_bo at 1.
            unfold ok_semstate.
            unfold bind at 3. unfold loc at 1. unfold bo at 1.
            unfold st at 1.
            unfold _get_bo at 1. unfold bind_s at 1. unfold bind at 3.
            unfold bind at 2.
            unfold bind at 2. unfold _get_bo at 1. unfold bind_s at 1.
            unfold bind at 2. unfold _get_bo at 1. unfold bind_s at 1.
            unfold _set_bo at 1. unfold ok_semstate.
            unfold bind at 2.
            unfold bind at 1. unfold loc. unfold bo. unfold st. simpl.
            simpl. rewrite same_bool.
            (* get the same projection relation as the one in hypothesis *)
            exact psrel.
          (* ConditionPassed(&proc->cpsr, cond) evaluates to false *)
          (* Skip statement from m7 to mfin, m7 = mfin *)
          inv main_p.
          (* expand ADC_step *)
          unfold S.ADC_step; unfold _get_st; unfold bind_s; unfold bind; simpl.
          rewrite cp_b; simpl.
          (* get the same projection relation as the one in hypothesis *)
          exact psrel.
Qed.

